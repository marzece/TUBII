/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from fifo_bettert.xcd on Fri Oct 20 11:53:28 1995 */
/* PART 3064PC84-125 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module fifo_ctrl
(SDOUT, SDIN, M2, RESET_n, BXREG_WR_n, BXREG_RD_n, BXREG_ADD, BWRITE_ENABLE_n, BWRITE_ADD_SEL_n, BREAD_ENABLE_n, BREAD_ADD_SEL_n, BMEM_WRITE_n, BMEM_READ_n, BD, BADD_OUT, P7, P8, P10, P11, PWRDWN_n, P28, P30, RDATA_n, RTRIG, P34, P36, P38, P44, P46, P48, P52, P53, PROGRAM_n, CCLK, P75, P76, P78);
   output SDOUT;
   input SDIN;
   output M2;
   input RESET_n;
   input BXREG_WR_n;
   input BXREG_RD_n;
   input [1:0] BXREG_ADD;
   output BWRITE_ENABLE_n;
   input BWRITE_ADD_SEL_n;
   output BREAD_ENABLE_n;
   input BREAD_ADD_SEL_n;
   input BMEM_WRITE_n;
   input BMEM_READ_n;
   inout [19:0] BD;
   inout [19:0] BADD_OUT;
   inout P7;
   inout P8;
   inout P10;
   inout P11;
   input PWRDWN_n;
   inout P28;
   inout P30;
   output RDATA_n;
   input RTRIG;
   inout P34;
   inout P36;
   inout P38;
   inout P44;
   inout P46;
   inout P48;
   inout P52;
   inout P53;
   input PROGRAM_n;
   input CCLK;
   inout P75;
   inout P76;
   inout P78;
wire [0:0] N125P_1_I93_1_I44_1_TQ;
wire [0:0] N125P_1_I93_1_I44_1_MD;
wire [0:0] N125P_1_I93_1_I44_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I44_1_I8_1_M0;
wire [0:0] N125P_1_I93_1_I43_1_TQ;
wire [0:0] N125P_1_I93_1_I43_1_MD;
wire [0:0] N125P_1_I93_1_I43_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I43_1_I8_1_M0;
wire [0:0] N125P_1_I93_1_I39_1_TQ;
wire [0:0] N125P_1_I93_1_I39_1_MD;
wire [0:0] N125P_1_I93_1_I39_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I39_1_I8_1_M0;
wire [0:0] N125P_1_I93_1_I36_1_TQ;
wire [0:0] N125P_1_I93_1_I36_1_MD;
wire [0:0] N125P_1_I93_1_I36_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I36_1_I8_1_M0;
wire [0:0] N125P_1_I93_1_I35_1_TQ;
wire [0:0] N125P_1_I93_1_I35_1_MD;
wire [0:0] N125P_1_I93_1_I35_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I35_1_I8_1_M0;
wire [0:0] N125P_1_I93_1_I31_1_TQ;
wire [0:0] N125P_1_I93_1_I31_1_MD;
wire [0:0] N125P_1_I93_1_I31_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I31_1_I8_1_M0;
wire [0:0] N125P_1_I93_1_I26_1_TQ;
wire [0:0] N125P_1_I93_1_I26_1_MD;
wire [0:0] N125P_1_I93_1_I26_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I26_1_I8_1_M0;
wire [0:0] N125P_1_I93_1_I25_1_TQ;
wire [0:0] N125P_1_I93_1_I25_1_MD;
wire [0:0] N125P_1_I93_1_I25_1_I8_1_M1;
wire [0:0] N125P_1_I93_1_I25_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I44_1_TQ;
wire [0:0] N125P_1_I92_1_I44_1_MD;
wire [0:0] N125P_1_I92_1_I44_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I44_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I43_1_TQ;
wire [0:0] N125P_1_I92_1_I43_1_MD;
wire [0:0] N125P_1_I92_1_I43_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I43_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I39_1_TQ;
wire [0:0] N125P_1_I92_1_I39_1_MD;
wire [0:0] N125P_1_I92_1_I39_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I39_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I36_1_TQ;
wire [0:0] N125P_1_I92_1_I36_1_MD;
wire [0:0] N125P_1_I92_1_I36_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I36_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I35_1_TQ;
wire [0:0] N125P_1_I92_1_I35_1_MD;
wire [0:0] N125P_1_I92_1_I35_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I35_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I31_1_TQ;
wire [0:0] N125P_1_I92_1_I31_1_MD;
wire [0:0] N125P_1_I92_1_I31_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I31_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I26_1_TQ;
wire [0:0] N125P_1_I92_1_I26_1_MD;
wire [0:0] N125P_1_I92_1_I26_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I26_1_I8_1_M0;
wire [0:0] N125P_1_I92_1_I25_1_TQ;
wire [0:0] N125P_1_I92_1_I25_1_MD;
wire [0:0] N125P_1_I92_1_I25_1_I8_1_M1;
wire [0:0] N125P_1_I92_1_I25_1_I8_1_M0;
wire [0:0] N125P_1_I90_1_I23_1_TQ;
wire [0:0] N125P_1_I90_1_I23_1_MD;
wire [0:0] N125P_1_I90_1_I23_1_I8_1_M1;
wire [0:0] N125P_1_I90_1_I23_1_I8_1_M0;
wire [0:0] N125P_1_I90_1_I22_1_TQ;
wire [0:0] N125P_1_I90_1_I22_1_MD;
wire [0:0] N125P_1_I90_1_I22_1_I8_1_M1;
wire [0:0] N125P_1_I90_1_I22_1_I8_1_M0;
wire [0:0] N125P_1_I90_1_I20_1_TQ;
wire [0:0] N125P_1_I90_1_I20_1_MD;
wire [0:0] N125P_1_I90_1_I20_1_I8_1_M1;
wire [0:0] N125P_1_I90_1_I20_1_I8_1_M0;
wire [0:0] N125P_1_I90_1_I18_1_TQ;
wire [0:0] N125P_1_I90_1_I18_1_MD;
wire [0:0] N125P_1_I90_1_I18_1_I8_1_M1;
wire [0:0] N125P_1_I90_1_I18_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I57_1_M1;
wire [0:0] N107P_1_108P_1_I57_1_M0;
wire [0:0] N107P_1_108P_1_I56_1_M1;
wire [0:0] N107P_1_108P_1_I56_1_M0;
wire [0:0] N107P_1_108P_1_I49_1_TQ;
wire [0:0] N107P_1_108P_1_I49_1_MD;
wire [0:0] N107P_1_108P_1_I49_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I49_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I46_1_TQ;
wire [0:0] N107P_1_108P_1_I46_1_MD;
wire [0:0] N107P_1_108P_1_I46_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I46_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I44_1_M1;
wire [0:0] N107P_1_108P_1_I44_1_M0;
wire [0:0] N107P_1_108P_1_I43_1_TQ;
wire [0:0] N107P_1_108P_1_I43_1_MD;
wire [0:0] N107P_1_108P_1_I43_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I43_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I42_1_TQ;
wire [0:0] N107P_1_108P_1_I42_1_MD;
wire [0:0] N107P_1_108P_1_I42_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I42_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I41_1_M1;
wire [0:0] N107P_1_108P_1_I41_1_M0;
wire [0:0] N107P_1_108P_1_I40_1_M1;
wire [0:0] N107P_1_108P_1_I40_1_M0;
wire [0:0] N107P_1_108P_1_I36_1_M1;
wire [0:0] N107P_1_108P_1_I36_1_M0;
wire [0:0] N107P_1_108P_1_I35_1_TQ;
wire [0:0] N107P_1_108P_1_I35_1_MD;
wire [0:0] N107P_1_108P_1_I35_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I35_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I34_1_TQ;
wire [0:0] N107P_1_108P_1_I34_1_MD;
wire [0:0] N107P_1_108P_1_I34_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I34_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I31_1_TQ;
wire [0:0] N107P_1_108P_1_I31_1_MD;
wire [0:0] N107P_1_108P_1_I31_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I31_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I30_1_M1;
wire [0:0] N107P_1_108P_1_I30_1_M0;
wire [0:0] N107P_1_108P_1_I29_1_TQ;
wire [0:0] N107P_1_108P_1_I29_1_MD;
wire [0:0] N107P_1_108P_1_I29_1_I8_1_M1;
wire [0:0] N107P_1_108P_1_I29_1_I8_1_M0;
wire [0:0] N107P_1_108P_1_I27_1_M1;
wire [0:0] N107P_1_108P_1_I27_1_M0;
wire [7:0] N107P_1_108P_1_D;
wire [0:0] N107P_1_107P_1_I57_1_M1;
wire [0:0] N107P_1_107P_1_I57_1_M0;
wire [0:0] N107P_1_107P_1_I56_1_M1;
wire [0:0] N107P_1_107P_1_I56_1_M0;
wire [0:0] N107P_1_107P_1_I49_1_TQ;
wire [0:0] N107P_1_107P_1_I49_1_MD;
wire [0:0] N107P_1_107P_1_I49_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I49_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I46_1_TQ;
wire [0:0] N107P_1_107P_1_I46_1_MD;
wire [0:0] N107P_1_107P_1_I46_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I46_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I44_1_M1;
wire [0:0] N107P_1_107P_1_I44_1_M0;
wire [0:0] N107P_1_107P_1_I43_1_TQ;
wire [0:0] N107P_1_107P_1_I43_1_MD;
wire [0:0] N107P_1_107P_1_I43_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I43_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I42_1_TQ;
wire [0:0] N107P_1_107P_1_I42_1_MD;
wire [0:0] N107P_1_107P_1_I42_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I42_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I41_1_M1;
wire [0:0] N107P_1_107P_1_I41_1_M0;
wire [0:0] N107P_1_107P_1_I40_1_M1;
wire [0:0] N107P_1_107P_1_I40_1_M0;
wire [0:0] N107P_1_107P_1_I36_1_M1;
wire [0:0] N107P_1_107P_1_I36_1_M0;
wire [0:0] N107P_1_107P_1_I35_1_TQ;
wire [0:0] N107P_1_107P_1_I35_1_MD;
wire [0:0] N107P_1_107P_1_I35_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I35_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I34_1_TQ;
wire [0:0] N107P_1_107P_1_I34_1_MD;
wire [0:0] N107P_1_107P_1_I34_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I34_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I31_1_TQ;
wire [0:0] N107P_1_107P_1_I31_1_MD;
wire [0:0] N107P_1_107P_1_I31_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I31_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I30_1_M1;
wire [0:0] N107P_1_107P_1_I30_1_M0;
wire [0:0] N107P_1_107P_1_I29_1_TQ;
wire [0:0] N107P_1_107P_1_I29_1_MD;
wire [0:0] N107P_1_107P_1_I29_1_I8_1_M1;
wire [0:0] N107P_1_107P_1_I29_1_I8_1_M0;
wire [0:0] N107P_1_107P_1_I27_1_M1;
wire [0:0] N107P_1_107P_1_I27_1_M0;
wire [7:0] N107P_1_107P_1_D;
wire [0:0] N107P_1_100P_1_I29_1_M1;
wire [0:0] N107P_1_100P_1_I29_1_M0;
wire [0:0] N107P_1_100P_1_I27_1_M1;
wire [0:0] N107P_1_100P_1_I27_1_M0;
wire [0:0] N107P_1_100P_1_I26_1_TQ;
wire [0:0] N107P_1_100P_1_I26_1_MD;
wire [0:0] N107P_1_100P_1_I26_1_I8_1_M1;
wire [0:0] N107P_1_100P_1_I26_1_I8_1_M0;
wire [0:0] N107P_1_100P_1_I25_1_TQ;
wire [0:0] N107P_1_100P_1_I25_1_MD;
wire [0:0] N107P_1_100P_1_I25_1_I8_1_M1;
wire [0:0] N107P_1_100P_1_I25_1_I8_1_M0;
wire [0:0] N107P_1_100P_1_I24_1_M1;
wire [0:0] N107P_1_100P_1_I24_1_M0;
wire [0:0] N107P_1_100P_1_I23_1_M1;
wire [0:0] N107P_1_100P_1_I23_1_M0;
wire [0:0] N107P_1_100P_1_I22_1_TQ;
wire [0:0] N107P_1_100P_1_I22_1_MD;
wire [0:0] N107P_1_100P_1_I22_1_I8_1_M1;
wire [0:0] N107P_1_100P_1_I22_1_I8_1_M0;
wire [0:0] N107P_1_100P_1_I18_1_TQ;
wire [0:0] N107P_1_100P_1_I18_1_MD;
wire [0:0] N107P_1_100P_1_I18_1_I8_1_M1;
wire [0:0] N107P_1_100P_1_I18_1_I8_1_M0;
wire [19:0] N107P_1_POINTER_ADDRESS;
wire [0:0] N91P_1_I93_1_I44_1_TQ;
wire [0:0] N91P_1_I93_1_I44_1_MD;
wire [0:0] N91P_1_I93_1_I44_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I44_1_I8_1_M0;
wire [0:0] N91P_1_I93_1_I43_1_TQ;
wire [0:0] N91P_1_I93_1_I43_1_MD;
wire [0:0] N91P_1_I93_1_I43_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I43_1_I8_1_M0;
wire [0:0] N91P_1_I93_1_I39_1_TQ;
wire [0:0] N91P_1_I93_1_I39_1_MD;
wire [0:0] N91P_1_I93_1_I39_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I39_1_I8_1_M0;
wire [0:0] N91P_1_I93_1_I36_1_TQ;
wire [0:0] N91P_1_I93_1_I36_1_MD;
wire [0:0] N91P_1_I93_1_I36_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I36_1_I8_1_M0;
wire [0:0] N91P_1_I93_1_I35_1_TQ;
wire [0:0] N91P_1_I93_1_I35_1_MD;
wire [0:0] N91P_1_I93_1_I35_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I35_1_I8_1_M0;
wire [0:0] N91P_1_I93_1_I31_1_TQ;
wire [0:0] N91P_1_I93_1_I31_1_MD;
wire [0:0] N91P_1_I93_1_I31_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I31_1_I8_1_M0;
wire [0:0] N91P_1_I93_1_I26_1_TQ;
wire [0:0] N91P_1_I93_1_I26_1_MD;
wire [0:0] N91P_1_I93_1_I26_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I26_1_I8_1_M0;
wire [0:0] N91P_1_I93_1_I25_1_TQ;
wire [0:0] N91P_1_I93_1_I25_1_MD;
wire [0:0] N91P_1_I93_1_I25_1_I8_1_M1;
wire [0:0] N91P_1_I93_1_I25_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I44_1_TQ;
wire [0:0] N91P_1_I92_1_I44_1_MD;
wire [0:0] N91P_1_I92_1_I44_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I44_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I43_1_TQ;
wire [0:0] N91P_1_I92_1_I43_1_MD;
wire [0:0] N91P_1_I92_1_I43_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I43_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I39_1_TQ;
wire [0:0] N91P_1_I92_1_I39_1_MD;
wire [0:0] N91P_1_I92_1_I39_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I39_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I36_1_TQ;
wire [0:0] N91P_1_I92_1_I36_1_MD;
wire [0:0] N91P_1_I92_1_I36_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I36_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I35_1_TQ;
wire [0:0] N91P_1_I92_1_I35_1_MD;
wire [0:0] N91P_1_I92_1_I35_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I35_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I31_1_TQ;
wire [0:0] N91P_1_I92_1_I31_1_MD;
wire [0:0] N91P_1_I92_1_I31_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I31_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I26_1_TQ;
wire [0:0] N91P_1_I92_1_I26_1_MD;
wire [0:0] N91P_1_I92_1_I26_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I26_1_I8_1_M0;
wire [0:0] N91P_1_I92_1_I25_1_TQ;
wire [0:0] N91P_1_I92_1_I25_1_MD;
wire [0:0] N91P_1_I92_1_I25_1_I8_1_M1;
wire [0:0] N91P_1_I92_1_I25_1_I8_1_M0;
wire [0:0] N91P_1_I90_1_I23_1_TQ;
wire [0:0] N91P_1_I90_1_I23_1_MD;
wire [0:0] N91P_1_I90_1_I23_1_I8_1_M1;
wire [0:0] N91P_1_I90_1_I23_1_I8_1_M0;
wire [0:0] N91P_1_I90_1_I22_1_TQ;
wire [0:0] N91P_1_I90_1_I22_1_MD;
wire [0:0] N91P_1_I90_1_I22_1_I8_1_M1;
wire [0:0] N91P_1_I90_1_I22_1_I8_1_M0;
wire [0:0] N91P_1_I90_1_I20_1_TQ;
wire [0:0] N91P_1_I90_1_I20_1_MD;
wire [0:0] N91P_1_I90_1_I20_1_I8_1_M1;
wire [0:0] N91P_1_I90_1_I20_1_I8_1_M0;
wire [0:0] N91P_1_I90_1_I18_1_TQ;
wire [0:0] N91P_1_I90_1_I18_1_MD;
wire [0:0] N91P_1_I90_1_I18_1_I8_1_M1;
wire [0:0] N91P_1_I90_1_I18_1_I8_1_M0;
wire [19:0] N73P_1_3P_1_M1;
wire [19:0] N73P_1_3P_1_M0;
wire [19:0] N73P_1_ADDRESS_OUT;
wire [0:0] N62P_1_16P_1_D3;
wire [0:0] N62P_1_16P_1_D2;
wire [0:0] N62P_1_1P_1_D3;
wire [1:0] XREG_ADD;
wire [19:0] XDT;
wire [19:0] WRITE_ADD;
wire [4:0] REG_CNTROL;
wire [19:0] READ_ADD;
wire [19:0] ADD_IN;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/peter/xilinx/fifo/fifo_ctrl/verilog_lib/fifo_ctrl.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

or2 N73P_1_3P_1_I5_1_20 (.o(N73P_1_ADDRESS_OUT[19]), .i0(N73P_1_3P_1_M1[19]), .i1(N73P_1_3P_1_M0[19]));
or2 N73P_1_3P_1_I5_1_19 (.i1(N73P_1_3P_1_M0[18]), .i0(N73P_1_3P_1_M1[18]), .o(N73P_1_ADDRESS_OUT[18]));
or2 N73P_1_3P_1_I5_1_18 (.i1(N73P_1_3P_1_M0[17]), .i0(N73P_1_3P_1_M1[17]), .o(N73P_1_ADDRESS_OUT[17]));
or2 N73P_1_3P_1_I5_1_17 (.i1(N73P_1_3P_1_M0[16]), .i0(N73P_1_3P_1_M1[16]), .o(N73P_1_ADDRESS_OUT[16]));
or2 N73P_1_3P_1_I5_1_16 (.i1(N73P_1_3P_1_M0[15]), .i0(N73P_1_3P_1_M1[15]), .o(N73P_1_ADDRESS_OUT[15]));
or2 N73P_1_3P_1_I5_1_15 (.i1(N73P_1_3P_1_M0[14]), .i0(N73P_1_3P_1_M1[14]), .o(N73P_1_ADDRESS_OUT[14]));
or2 N73P_1_3P_1_I5_1_14 (.i1(N73P_1_3P_1_M0[13]), .i0(N73P_1_3P_1_M1[13]), .o(N73P_1_ADDRESS_OUT[13]));
or2 N73P_1_3P_1_I5_1_13 (.i1(N73P_1_3P_1_M0[12]), .i0(N73P_1_3P_1_M1[12]), .o(N73P_1_ADDRESS_OUT[12]));
or2 N73P_1_3P_1_I5_1_12 (.i1(N73P_1_3P_1_M0[11]), .i0(N73P_1_3P_1_M1[11]), .o(N73P_1_ADDRESS_OUT[11]));
or2 N73P_1_3P_1_I5_1_11 (.i1(N73P_1_3P_1_M0[10]), .i0(N73P_1_3P_1_M1[10]), .o(N73P_1_ADDRESS_OUT[10]));
or2 N73P_1_3P_1_I5_1_10 (.i1(N73P_1_3P_1_M0[9]), .i0(N73P_1_3P_1_M1[9]), .o(N73P_1_ADDRESS_OUT[9]));
or2 N73P_1_3P_1_I5_1_9 (.i1(N73P_1_3P_1_M0[8]), .i0(N73P_1_3P_1_M1[8]), .o(N73P_1_ADDRESS_OUT[8]));
or2 N73P_1_3P_1_I5_1_8 (.i1(N73P_1_3P_1_M0[7]), .i0(N73P_1_3P_1_M1[7]), .o(N73P_1_ADDRESS_OUT[7]));
or2 N73P_1_3P_1_I5_1_7 (.i1(N73P_1_3P_1_M0[6]), .i0(N73P_1_3P_1_M1[6]), .o(N73P_1_ADDRESS_OUT[6]));
or2 N73P_1_3P_1_I5_1_6 (.i1(N73P_1_3P_1_M0[5]), .i0(N73P_1_3P_1_M1[5]), .o(N73P_1_ADDRESS_OUT[5]));
or2 N73P_1_3P_1_I5_1_5 (.i1(N73P_1_3P_1_M0[4]), .i0(N73P_1_3P_1_M1[4]), .o(N73P_1_ADDRESS_OUT[4]));
or2 N73P_1_3P_1_I5_1_4 (.i1(N73P_1_3P_1_M0[3]), .i0(N73P_1_3P_1_M1[3]), .o(N73P_1_ADDRESS_OUT[3]));
or2 N73P_1_3P_1_I5_1_3 (.i1(N73P_1_3P_1_M0[2]), .i0(N73P_1_3P_1_M1[2]), .o(N73P_1_ADDRESS_OUT[2]));
or2 N73P_1_3P_1_I5_1_2 (.i1(N73P_1_3P_1_M0[1]), .i0(N73P_1_3P_1_M1[1]), .o(N73P_1_ADDRESS_OUT[1]));
or2 N73P_1_3P_1_I5_1_1 (.i1(N73P_1_3P_1_M0[0]), .i0(N73P_1_3P_1_M1[0]), .o(N73P_1_ADDRESS_OUT[0]));
and2b1 N73P_1_3P_1_I7_1_20 (.o(N73P_1_3P_1_M0[19]), .i0(N_WRITE_ADD_SEL), .i1(WRITE_ADD[19]));
and2b1 N73P_1_3P_1_I7_1_19 (.i1(WRITE_ADD[18]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[18]));
and2b1 N73P_1_3P_1_I7_1_18 (.i1(WRITE_ADD[17]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[17]));
and2b1 N73P_1_3P_1_I7_1_17 (.i1(WRITE_ADD[16]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[16]));
and2b1 N73P_1_3P_1_I7_1_16 (.i1(WRITE_ADD[15]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[15]));
and2b1 N73P_1_3P_1_I7_1_15 (.i1(WRITE_ADD[14]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[14]));
and2b1 N73P_1_3P_1_I7_1_14 (.i1(WRITE_ADD[13]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[13]));
and2b1 N73P_1_3P_1_I7_1_13 (.i1(WRITE_ADD[12]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[12]));
and2b1 N73P_1_3P_1_I7_1_12 (.i1(WRITE_ADD[11]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[11]));
and2b1 N73P_1_3P_1_I7_1_11 (.i1(WRITE_ADD[10]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[10]));
and2b1 N73P_1_3P_1_I7_1_10 (.i1(WRITE_ADD[9]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[9]));
and2b1 N73P_1_3P_1_I7_1_9 (.i1(WRITE_ADD[8]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[8]));
and2b1 N73P_1_3P_1_I7_1_8 (.i1(WRITE_ADD[7]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[7]));
and2b1 N73P_1_3P_1_I7_1_7 (.i1(WRITE_ADD[6]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[6]));
and2b1 N73P_1_3P_1_I7_1_6 (.i1(WRITE_ADD[5]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[5]));
and2b1 N73P_1_3P_1_I7_1_5 (.i1(WRITE_ADD[4]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[4]));
and2b1 N73P_1_3P_1_I7_1_4 (.i1(WRITE_ADD[3]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[3]));
and2b1 N73P_1_3P_1_I7_1_3 (.i1(WRITE_ADD[2]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[2]));
and2b1 N73P_1_3P_1_I7_1_2 (.i1(WRITE_ADD[1]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[1]));
and2b1 N73P_1_3P_1_I7_1_1 (.i1(WRITE_ADD[0]), .i0(N_WRITE_ADD_SEL), .o(N73P_1_3P_1_M0[0]));
and2 N73P_1_3P_1_I6_1_20 (.o(N73P_1_3P_1_M1[19]), .i0(READ_ADD[19]), .i1(N_WRITE_ADD_SEL));
and2 N73P_1_3P_1_I6_1_19 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[18]), .o(N73P_1_3P_1_M1[18]));
and2 N73P_1_3P_1_I6_1_18 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[17]), .o(N73P_1_3P_1_M1[17]));
and2 N73P_1_3P_1_I6_1_17 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[16]), .o(N73P_1_3P_1_M1[16]));
and2 N73P_1_3P_1_I6_1_16 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[15]), .o(N73P_1_3P_1_M1[15]));
and2 N73P_1_3P_1_I6_1_15 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[14]), .o(N73P_1_3P_1_M1[14]));
and2 N73P_1_3P_1_I6_1_14 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[13]), .o(N73P_1_3P_1_M1[13]));
and2 N73P_1_3P_1_I6_1_13 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[12]), .o(N73P_1_3P_1_M1[12]));
and2 N73P_1_3P_1_I6_1_12 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[11]), .o(N73P_1_3P_1_M1[11]));
and2 N73P_1_3P_1_I6_1_11 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[10]), .o(N73P_1_3P_1_M1[10]));
and2 N73P_1_3P_1_I6_1_10 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[9]), .o(N73P_1_3P_1_M1[9]));
and2 N73P_1_3P_1_I6_1_9 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[8]), .o(N73P_1_3P_1_M1[8]));
and2 N73P_1_3P_1_I6_1_8 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[7]), .o(N73P_1_3P_1_M1[7]));
and2 N73P_1_3P_1_I6_1_7 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[6]), .o(N73P_1_3P_1_M1[6]));
and2 N73P_1_3P_1_I6_1_6 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[5]), .o(N73P_1_3P_1_M1[5]));
and2 N73P_1_3P_1_I6_1_5 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[4]), .o(N73P_1_3P_1_M1[4]));
and2 N73P_1_3P_1_I6_1_4 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[3]), .o(N73P_1_3P_1_M1[3]));
and2 N73P_1_3P_1_I6_1_3 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[2]), .o(N73P_1_3P_1_M1[2]));
and2 N73P_1_3P_1_I6_1_2 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[1]), .o(N73P_1_3P_1_M1[1]));
and2 N73P_1_3P_1_I6_1_1 (.i1(N_WRITE_ADD_SEL), .i0(READ_ADD[0]), .o(N73P_1_3P_1_M1[0]));
ibuf N73P_1_9P_1_20 (.i(BD[19]), .o(ADD_IN[19]));
ibuf N73P_1_9P_1_19 (.o(ADD_IN[18]), .i(BD[18]));
ibuf N73P_1_9P_1_18 (.o(ADD_IN[17]), .i(BD[17]));
ibuf N73P_1_9P_1_17 (.o(ADD_IN[16]), .i(BD[16]));
ibuf N73P_1_9P_1_16 (.o(ADD_IN[15]), .i(BD[15]));
ibuf N73P_1_9P_1_15 (.o(ADD_IN[14]), .i(BD[14]));
ibuf N73P_1_9P_1_14 (.o(ADD_IN[13]), .i(BD[13]));
ibuf N73P_1_9P_1_13 (.o(ADD_IN[12]), .i(BD[12]));
ibuf N73P_1_9P_1_12 (.o(ADD_IN[11]), .i(BD[11]));
ibuf N73P_1_9P_1_11 (.o(ADD_IN[10]), .i(BD[10]));
ibuf N73P_1_9P_1_10 (.o(ADD_IN[9]), .i(BD[9]));
ibuf N73P_1_9P_1_9 (.o(ADD_IN[8]), .i(BD[8]));
ibuf N73P_1_9P_1_8 (.o(ADD_IN[7]), .i(BD[7]));
ibuf N73P_1_9P_1_7 (.o(ADD_IN[6]), .i(BD[6]));
ibuf N73P_1_9P_1_6 (.o(ADD_IN[5]), .i(BD[5]));
ibuf N73P_1_9P_1_5 (.o(ADD_IN[4]), .i(BD[4]));
ibuf N73P_1_9P_1_4 (.o(ADD_IN[3]), .i(BD[3]));
ibuf N73P_1_9P_1_3 (.o(ADD_IN[2]), .i(BD[2]));
ibuf N73P_1_9P_1_2 (.o(ADD_IN[1]), .i(BD[1]));
ibuf N73P_1_9P_1_1 (.o(ADD_IN[0]), .i(BD[0]));
obuft N73P_1_30P_1_10 (.i(N73P_1_ADDRESS_OUT[9]), .o(BADD_OUT[9]), .t(N73P_1_N_ADD_OUT_ENABLE));
obuft N73P_1_30P_1_9 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[8]), .i(N73P_1_ADDRESS_OUT[8]));
obuft N73P_1_30P_1_8 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[7]), .i(N73P_1_ADDRESS_OUT[7]));
obuft N73P_1_30P_1_7 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[6]), .i(N73P_1_ADDRESS_OUT[6]));
obuft N73P_1_30P_1_6 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[5]), .i(N73P_1_ADDRESS_OUT[5]));
obuft N73P_1_30P_1_5 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[4]), .i(N73P_1_ADDRESS_OUT[4]));
obuft N73P_1_30P_1_4 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[3]), .i(N73P_1_ADDRESS_OUT[3]));
obuft N73P_1_30P_1_3 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[2]), .i(N73P_1_ADDRESS_OUT[2]));
obuft N73P_1_30P_1_2 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[1]), .i(N73P_1_ADDRESS_OUT[1]));
obuft N73P_1_30P_1_1 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[0]), .i(N73P_1_ADDRESS_OUT[0]));
obuft N73P_1_29P_1_10 (.i(N73P_1_ADDRESS_OUT[19]), .o(BADD_OUT[19]), .t(N73P_1_N_ADD_OUT_ENABLE));
obuft N73P_1_29P_1_9 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[18]), .i(N73P_1_ADDRESS_OUT[18]));
obuft N73P_1_29P_1_8 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[17]), .i(N73P_1_ADDRESS_OUT[17]));
obuft N73P_1_29P_1_7 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[16]), .i(N73P_1_ADDRESS_OUT[16]));
obuft N73P_1_29P_1_6 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[15]), .i(N73P_1_ADDRESS_OUT[15]));
obuft N73P_1_29P_1_5 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[14]), .i(N73P_1_ADDRESS_OUT[14]));
obuft N73P_1_29P_1_4 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[13]), .i(N73P_1_ADDRESS_OUT[13]));
obuft N73P_1_29P_1_3 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[12]), .i(N73P_1_ADDRESS_OUT[12]));
obuft N73P_1_29P_1_2 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[11]), .i(N73P_1_ADDRESS_OUT[11]));
obuft N73P_1_29P_1_1 (.t(N73P_1_N_ADD_OUT_ENABLE), .o(BADD_OUT[10]), .i(N73P_1_ADDRESS_OUT[10]));
obuft N73P_1_8P_1_20 (.i(XDT[19]), .o(BD[19]), .t(N_XREG_RD));
obuft N73P_1_8P_1_19 (.t(N_XREG_RD), .o(BD[18]), .i(XDT[18]));
obuft N73P_1_8P_1_18 (.t(N_XREG_RD), .o(BD[17]), .i(XDT[17]));
obuft N73P_1_8P_1_17 (.t(N_XREG_RD), .o(BD[16]), .i(XDT[16]));
obuft N73P_1_8P_1_16 (.t(N_XREG_RD), .o(BD[15]), .i(XDT[15]));
obuft N73P_1_8P_1_15 (.t(N_XREG_RD), .o(BD[14]), .i(XDT[14]));
obuft N73P_1_8P_1_14 (.t(N_XREG_RD), .o(BD[13]), .i(XDT[13]));
obuft N73P_1_8P_1_13 (.t(N_XREG_RD), .o(BD[12]), .i(XDT[12]));
obuft N73P_1_8P_1_12 (.t(N_XREG_RD), .o(BD[11]), .i(XDT[11]));
obuft N73P_1_8P_1_11 (.t(N_XREG_RD), .o(BD[10]), .i(XDT[10]));
obuft N73P_1_8P_1_10 (.t(N_XREG_RD), .o(BD[9]), .i(XDT[9]));
obuft N73P_1_8P_1_9 (.t(N_XREG_RD), .o(BD[8]), .i(XDT[8]));
obuft N73P_1_8P_1_8 (.t(N_XREG_RD), .o(BD[7]), .i(XDT[7]));
obuft N73P_1_8P_1_7 (.t(N_XREG_RD), .o(BD[6]), .i(XDT[6]));
obuft N73P_1_8P_1_6 (.t(N_XREG_RD), .o(BD[5]), .i(XDT[5]));
obuft N73P_1_8P_1_5 (.t(N_XREG_RD), .o(BD[4]), .i(XDT[4]));
obuft N73P_1_8P_1_4 (.t(N_XREG_RD), .o(BD[3]), .i(XDT[3]));
obuft N73P_1_8P_1_3 (.t(N_XREG_RD), .o(BD[2]), .i(XDT[2]));
obuft N73P_1_8P_1_2 (.t(N_XREG_RD), .o(BD[1]), .i(XDT[1]));
obuft N73P_1_8P_1_1 (.t(N_XREG_RD), .o(BD[0]), .i(XDT[0]));
and2b1 N73P_1_25P_1 (.o(N73P_1_UN_1_AND2B1_25P_O), .i0(N_READ_ADD_SEL), .i1(WRITE_ENABLE));
and2b1 N73P_1_26P_1 (.o(N73P_1_UN_1_AND2B1_26P_O), .i0(N_WRITE_ADD_SEL), .i1(READ_ENABLE));
nor2 N73P_1_20P_1 (.o(N73P_1_N_ADD_OUT_ENABLE), .i0(N73P_1_UN_1_AND2B1_26P_O), .i1(N73P_1_UN_1_AND2B1_25P_O));
and3b1 N62P_1_16P_1_I13_1 (.i2(N62P_1_UN_1_D2_4E_16P_E), .o(N62P_1_UN_1_D2_4E_16P_D1), .i0(XREG_ADD[1]), .i1(XREG_ADD[0]));
and3b1 N62P_1_16P_1_I12_1 (.i2(N62P_1_UN_1_D2_4E_16P_E), .o(N62P_1_16P_1_D2[0]), .i0(XREG_ADD[0]), .i1(XREG_ADD[1]));
and3b2 N62P_1_16P_1_I9_1 (.i2(N62P_1_UN_1_D2_4E_16P_E), .o(N62P_1_UN_1_D2_4E_16P_D0), .i1(XREG_ADD[0]), .i0(XREG_ADD[1]));
and3 N62P_1_16P_1_I11_1 (.i2(N62P_1_UN_1_D2_4E_16P_E), .o(N62P_1_16P_1_D3[0]), .i0(XREG_ADD[1]), .i1(XREG_ADD[0]));
and3b1 N62P_1_1P_1_I13_1 (.i2(N62P_1_UN_1_D2_4E_1P_E), .o(N62P_1_UN_1_D2_4E_1P_D1), .i0(XREG_ADD[1]), .i1(XREG_ADD[0]));
and3b1 N62P_1_1P_1_I12_1 (.i2(N62P_1_UN_1_D2_4E_1P_E), .o(N62P_1_UN_1_D2_4E_1P_D2), .i0(XREG_ADD[0]), .i1(XREG_ADD[1]));
and3b2 N62P_1_1P_1_I9_1 (.i2(N62P_1_UN_1_D2_4E_1P_E), .o(N62P_1_UN_1_D2_4E_1P_D0), .i1(XREG_ADD[0]), .i0(XREG_ADD[1]));
and3 N62P_1_1P_1_I11_1 (.i2(N62P_1_UN_1_D2_4E_1P_E), .o(N62P_1_1P_1_D3[0]), .i0(XREG_ADD[1]), .i1(XREG_ADD[0]));
inv N62P_1_31P_1 (.i(N62P_1_UN_1_D2_4E_16P_D1), .o(REG_CNTROL[3]));
inv N62P_1_30P_1 (.i(N62P_1_UN_1_D2_4E_16P_D0), .o(REG_CNTROL[4]));
inv N62P_1_29P_1 (.i(N62P_1_UN_1_D2_4E_1P_D2), .o(REG_CNTROL[2]));
inv N62P_1_28P_1 (.i(N62P_1_UN_1_D2_4E_1P_D1), .o(REG_CNTROL[0]));
inv N62P_1_27P_1 (.i(N62P_1_UN_1_D2_4E_1P_D0), .o(REG_CNTROL[1]));
inv N62P_1_33P_1 (.i(N_XREG_WR), .o(N62P_1_UN_1_D2_4E_16P_E));
inv N62P_1_32P_1 (.i(N_XREG_RD), .o(N62P_1_UN_1_D2_4E_1P_E));
or2 N91P_1_I93_1_I44_1_I8_1_I5_1 (.o(N91P_1_I93_1_I44_1_MD[0]), .i0(N91P_1_I93_1_I44_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I44_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I44_1_I8_1_I7_1 (.o(N91P_1_I93_1_I44_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I44_1_TQ[0]));
and2 N91P_1_I93_1_I44_1_I8_1_I6_1 (.o(N91P_1_I93_1_I44_1_I8_1_M1[0]), .i0(ADD_IN[14]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I44_1_I12_1 (.q(READ_ADD[14]), .d(N91P_1_I93_1_I44_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I44_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I44_1_I13_1 (.o(N91P_1_I93_1_I44_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I44_1_I9_1 (.o(N91P_1_I93_1_I44_1_TQ[0]), .i0(N91P_1_I93_1_T6), .i1(READ_ADD[14]));
or2 N91P_1_I93_1_I43_1_I8_1_I5_1 (.o(N91P_1_I93_1_I43_1_MD[0]), .i0(N91P_1_I93_1_I43_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I43_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I43_1_I8_1_I7_1 (.o(N91P_1_I93_1_I43_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I43_1_TQ[0]));
and2 N91P_1_I93_1_I43_1_I8_1_I6_1 (.o(N91P_1_I93_1_I43_1_I8_1_M1[0]), .i0(ADD_IN[13]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I43_1_I12_1 (.q(READ_ADD[13]), .d(N91P_1_I93_1_I43_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I43_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I43_1_I13_1 (.o(N91P_1_I93_1_I43_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I43_1_I9_1 (.o(N91P_1_I93_1_I43_1_TQ[0]), .i0(N91P_1_I93_1_T5), .i1(READ_ADD[13]));
or2 N91P_1_I93_1_I39_1_I8_1_I5_1 (.o(N91P_1_I93_1_I39_1_MD[0]), .i0(N91P_1_I93_1_I39_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I39_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I39_1_I8_1_I7_1 (.o(N91P_1_I93_1_I39_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I39_1_TQ[0]));
and2 N91P_1_I93_1_I39_1_I8_1_I6_1 (.o(N91P_1_I93_1_I39_1_I8_1_M1[0]), .i0(ADD_IN[15]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I39_1_I12_1 (.q(READ_ADD[15]), .d(N91P_1_I93_1_I39_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I39_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I39_1_I13_1 (.o(N91P_1_I93_1_I39_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I39_1_I9_1 (.o(N91P_1_I93_1_I39_1_TQ[0]), .i0(N91P_1_I93_1_T7), .i1(READ_ADD[15]));
or2 N91P_1_I93_1_I36_1_I8_1_I5_1 (.o(N91P_1_I93_1_I36_1_MD[0]), .i0(N91P_1_I93_1_I36_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I36_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I36_1_I8_1_I7_1 (.o(N91P_1_I93_1_I36_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I36_1_TQ[0]));
and2 N91P_1_I93_1_I36_1_I8_1_I6_1 (.o(N91P_1_I93_1_I36_1_I8_1_M1[0]), .i0(ADD_IN[11]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I36_1_I12_1 (.q(READ_ADD[11]), .d(N91P_1_I93_1_I36_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I36_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I36_1_I13_1 (.o(N91P_1_I93_1_I36_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I36_1_I9_1 (.o(N91P_1_I93_1_I36_1_TQ[0]), .i0(N91P_1_I93_1_T3), .i1(READ_ADD[11]));
or2 N91P_1_I93_1_I35_1_I8_1_I5_1 (.o(N91P_1_I93_1_I35_1_MD[0]), .i0(N91P_1_I93_1_I35_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I35_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I35_1_I8_1_I7_1 (.o(N91P_1_I93_1_I35_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I35_1_TQ[0]));
and2 N91P_1_I93_1_I35_1_I8_1_I6_1 (.o(N91P_1_I93_1_I35_1_I8_1_M1[0]), .i0(ADD_IN[8]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I35_1_I12_1 (.q(READ_ADD[8]), .d(N91P_1_I93_1_I35_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I35_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I35_1_I13_1 (.o(N91P_1_I93_1_I35_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I35_1_I9_1 (.o(N91P_1_I93_1_I35_1_TQ[0]), .i0(XVDD), .i1(READ_ADD[8]));
or2 N91P_1_I93_1_I31_1_I8_1_I5_1 (.o(N91P_1_I93_1_I31_1_MD[0]), .i0(N91P_1_I93_1_I31_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I31_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I31_1_I8_1_I7_1 (.o(N91P_1_I93_1_I31_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I31_1_TQ[0]));
and2 N91P_1_I93_1_I31_1_I8_1_I6_1 (.o(N91P_1_I93_1_I31_1_I8_1_M1[0]), .i0(ADD_IN[9]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I31_1_I12_1 (.q(READ_ADD[9]), .d(N91P_1_I93_1_I31_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I31_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I31_1_I13_1 (.o(N91P_1_I93_1_I31_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I31_1_I9_1 (.o(N91P_1_I93_1_I31_1_TQ[0]), .i0(READ_ADD[8]), .i1(READ_ADD[9]));
or2 N91P_1_I93_1_I26_1_I8_1_I5_1 (.o(N91P_1_I93_1_I26_1_MD[0]), .i0(N91P_1_I93_1_I26_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I26_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I26_1_I8_1_I7_1 (.o(N91P_1_I93_1_I26_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I26_1_TQ[0]));
and2 N91P_1_I93_1_I26_1_I8_1_I6_1 (.o(N91P_1_I93_1_I26_1_I8_1_M1[0]), .i0(ADD_IN[10]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I26_1_I12_1 (.q(READ_ADD[10]), .d(N91P_1_I93_1_I26_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I26_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I26_1_I13_1 (.o(N91P_1_I93_1_I26_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I26_1_I9_1 (.o(N91P_1_I93_1_I26_1_TQ[0]), .i0(N91P_1_I93_1_T2), .i1(READ_ADD[10]));
or2 N91P_1_I93_1_I25_1_I8_1_I5_1 (.o(N91P_1_I93_1_I25_1_MD[0]), .i0(N91P_1_I93_1_I25_1_I8_1_M1[0]), .i1(N91P_1_I93_1_I25_1_I8_1_M0[0]));
and2b1 N91P_1_I93_1_I25_1_I8_1_I7_1 (.o(N91P_1_I93_1_I25_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I93_1_I25_1_TQ[0]));
and2 N91P_1_I93_1_I25_1_I8_1_I6_1 (.o(N91P_1_I93_1_I25_1_I8_1_M1[0]), .i0(ADD_IN[12]), .i1(N91P_1_LD));
fdce N91P_1_I93_1_I25_1_I12_1 (.q(READ_ADD[12]), .d(N91P_1_I93_1_I25_1_MD[0]), .c(READ_CU), .ce(N91P_1_I93_1_I25_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I93_1_I25_1_I13_1 (.o(N91P_1_I93_1_I25_1_L_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_LD));
xor2 N91P_1_I93_1_I25_1_I9_1 (.o(N91P_1_I93_1_I25_1_TQ[0]), .i0(N91P_1_I93_1_T4), .i1(READ_ADD[12]));
and3 N91P_1_I93_1_I29_1 (.i2(READ_ADD[8]), .o(N91P_1_I93_1_T3), .i0(READ_ADD[10]), .i1(READ_ADD[9]));
and3 N91P_1_I93_1_I27_1 (.i2(N91P_1_I93_1_T4), .o(N91P_1_I93_1_T6), .i0(READ_ADD[13]), .i1(READ_ADD[12]));
and4 N91P_1_I93_1_I38_1 (.i2(READ_ADD[9]), .i3(READ_ADD[8]), .o(N91P_1_I93_1_T4), .i0(READ_ADD[11]), .i1(READ_ADD[10]));
and4 N91P_1_I93_1_I33_1 (.i2(READ_ADD[12]), .i3(N91P_1_I93_1_T4), .o(N91P_1_I93_1_T7), .i0(READ_ADD[14]), .i1(READ_ADD[13]));
and5 N91P_1_I93_1_I37_1 (.i4(N91P_1_I93_1_T4), .i2(READ_ADD[13]), .i3(READ_ADD[12]), .o(N91P_1_I93_1_TC), .i0(READ_ADD[15]), .i1(READ_ADD[14]));
and2 N91P_1_I93_1_I34_1 (.o(N91P_1_I93_1_T5), .i0(READ_ADD[12]), .i1(N91P_1_I93_1_T4));
and2 N91P_1_I93_1_I32_1 (.o(N91P_1_UN_1_CB4CLE_I90_CE), .i0(N91P_1_UN_1_CB8CLE_I92_CEO), .i1(N91P_1_I93_1_TC));
and2 N91P_1_I93_1_I30_1 (.o(N91P_1_I93_1_T2), .i0(READ_ADD[9]), .i1(READ_ADD[8]));
or2 N91P_1_I92_1_I44_1_I8_1_I5_1 (.o(N91P_1_I92_1_I44_1_MD[0]), .i0(N91P_1_I92_1_I44_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I44_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I44_1_I8_1_I7_1 (.o(N91P_1_I92_1_I44_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I44_1_TQ[0]));
and2 N91P_1_I92_1_I44_1_I8_1_I6_1 (.o(N91P_1_I92_1_I44_1_I8_1_M1[0]), .i0(ADD_IN[6]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I44_1_I12_1 (.q(READ_ADD[6]), .d(N91P_1_I92_1_I44_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I44_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I44_1_I13_1 (.o(N91P_1_I92_1_I44_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I44_1_I9_1 (.o(N91P_1_I92_1_I44_1_TQ[0]), .i0(N91P_1_I92_1_T6), .i1(READ_ADD[6]));
or2 N91P_1_I92_1_I43_1_I8_1_I5_1 (.o(N91P_1_I92_1_I43_1_MD[0]), .i0(N91P_1_I92_1_I43_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I43_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I43_1_I8_1_I7_1 (.o(N91P_1_I92_1_I43_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I43_1_TQ[0]));
and2 N91P_1_I92_1_I43_1_I8_1_I6_1 (.o(N91P_1_I92_1_I43_1_I8_1_M1[0]), .i0(ADD_IN[5]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I43_1_I12_1 (.q(READ_ADD[5]), .d(N91P_1_I92_1_I43_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I43_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I43_1_I13_1 (.o(N91P_1_I92_1_I43_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I43_1_I9_1 (.o(N91P_1_I92_1_I43_1_TQ[0]), .i0(N91P_1_I92_1_T5), .i1(READ_ADD[5]));
or2 N91P_1_I92_1_I39_1_I8_1_I5_1 (.o(N91P_1_I92_1_I39_1_MD[0]), .i0(N91P_1_I92_1_I39_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I39_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I39_1_I8_1_I7_1 (.o(N91P_1_I92_1_I39_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I39_1_TQ[0]));
and2 N91P_1_I92_1_I39_1_I8_1_I6_1 (.o(N91P_1_I92_1_I39_1_I8_1_M1[0]), .i0(ADD_IN[7]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I39_1_I12_1 (.q(READ_ADD[7]), .d(N91P_1_I92_1_I39_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I39_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I39_1_I13_1 (.o(N91P_1_I92_1_I39_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I39_1_I9_1 (.o(N91P_1_I92_1_I39_1_TQ[0]), .i0(N91P_1_I92_1_T7), .i1(READ_ADD[7]));
or2 N91P_1_I92_1_I36_1_I8_1_I5_1 (.o(N91P_1_I92_1_I36_1_MD[0]), .i0(N91P_1_I92_1_I36_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I36_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I36_1_I8_1_I7_1 (.o(N91P_1_I92_1_I36_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I36_1_TQ[0]));
and2 N91P_1_I92_1_I36_1_I8_1_I6_1 (.o(N91P_1_I92_1_I36_1_I8_1_M1[0]), .i0(ADD_IN[3]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I36_1_I12_1 (.q(READ_ADD[3]), .d(N91P_1_I92_1_I36_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I36_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I36_1_I13_1 (.o(N91P_1_I92_1_I36_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I36_1_I9_1 (.o(N91P_1_I92_1_I36_1_TQ[0]), .i0(N91P_1_I92_1_T3), .i1(READ_ADD[3]));
or2 N91P_1_I92_1_I35_1_I8_1_I5_1 (.o(N91P_1_I92_1_I35_1_MD[0]), .i0(N91P_1_I92_1_I35_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I35_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I35_1_I8_1_I7_1 (.o(N91P_1_I92_1_I35_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I35_1_TQ[0]));
and2 N91P_1_I92_1_I35_1_I8_1_I6_1 (.o(N91P_1_I92_1_I35_1_I8_1_M1[0]), .i0(ADD_IN[0]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I35_1_I12_1 (.q(READ_ADD[0]), .d(N91P_1_I92_1_I35_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I35_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I35_1_I13_1 (.o(N91P_1_I92_1_I35_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I35_1_I9_1 (.o(N91P_1_I92_1_I35_1_TQ[0]), .i0(XVDD), .i1(READ_ADD[0]));
or2 N91P_1_I92_1_I31_1_I8_1_I5_1 (.o(N91P_1_I92_1_I31_1_MD[0]), .i0(N91P_1_I92_1_I31_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I31_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I31_1_I8_1_I7_1 (.o(N91P_1_I92_1_I31_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I31_1_TQ[0]));
and2 N91P_1_I92_1_I31_1_I8_1_I6_1 (.o(N91P_1_I92_1_I31_1_I8_1_M1[0]), .i0(ADD_IN[1]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I31_1_I12_1 (.q(READ_ADD[1]), .d(N91P_1_I92_1_I31_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I31_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I31_1_I13_1 (.o(N91P_1_I92_1_I31_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I31_1_I9_1 (.o(N91P_1_I92_1_I31_1_TQ[0]), .i0(READ_ADD[0]), .i1(READ_ADD[1]));
or2 N91P_1_I92_1_I26_1_I8_1_I5_1 (.o(N91P_1_I92_1_I26_1_MD[0]), .i0(N91P_1_I92_1_I26_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I26_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I26_1_I8_1_I7_1 (.o(N91P_1_I92_1_I26_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I26_1_TQ[0]));
and2 N91P_1_I92_1_I26_1_I8_1_I6_1 (.o(N91P_1_I92_1_I26_1_I8_1_M1[0]), .i0(ADD_IN[2]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I26_1_I12_1 (.q(READ_ADD[2]), .d(N91P_1_I92_1_I26_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I26_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I26_1_I13_1 (.o(N91P_1_I92_1_I26_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I26_1_I9_1 (.o(N91P_1_I92_1_I26_1_TQ[0]), .i0(N91P_1_I92_1_T2), .i1(READ_ADD[2]));
or2 N91P_1_I92_1_I25_1_I8_1_I5_1 (.o(N91P_1_I92_1_I25_1_MD[0]), .i0(N91P_1_I92_1_I25_1_I8_1_M1[0]), .i1(N91P_1_I92_1_I25_1_I8_1_M0[0]));
and2b1 N91P_1_I92_1_I25_1_I8_1_I7_1 (.o(N91P_1_I92_1_I25_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I92_1_I25_1_TQ[0]));
and2 N91P_1_I92_1_I25_1_I8_1_I6_1 (.o(N91P_1_I92_1_I25_1_I8_1_M1[0]), .i0(ADD_IN[4]), .i1(N91P_1_LD));
fdce N91P_1_I92_1_I25_1_I12_1 (.q(READ_ADD[4]), .d(N91P_1_I92_1_I25_1_MD[0]), .c(READ_CU), .ce(N91P_1_I92_1_I25_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I92_1_I25_1_I13_1 (.o(N91P_1_I92_1_I25_1_L_CE), .i0(READ_ENABLE), .i1(N91P_1_LD));
xor2 N91P_1_I92_1_I25_1_I9_1 (.o(N91P_1_I92_1_I25_1_TQ[0]), .i0(N91P_1_I92_1_T4), .i1(READ_ADD[4]));
and3 N91P_1_I92_1_I29_1 (.i2(READ_ADD[0]), .o(N91P_1_I92_1_T3), .i0(READ_ADD[2]), .i1(READ_ADD[1]));
and3 N91P_1_I92_1_I27_1 (.i2(N91P_1_I92_1_T4), .o(N91P_1_I92_1_T6), .i0(READ_ADD[5]), .i1(READ_ADD[4]));
and4 N91P_1_I92_1_I38_1 (.i2(READ_ADD[1]), .i3(READ_ADD[0]), .o(N91P_1_I92_1_T4), .i0(READ_ADD[3]), .i1(READ_ADD[2]));
and4 N91P_1_I92_1_I33_1 (.i2(READ_ADD[4]), .i3(N91P_1_I92_1_T4), .o(N91P_1_I92_1_T7), .i0(READ_ADD[6]), .i1(READ_ADD[5]));
and5 N91P_1_I92_1_I37_1 (.i4(N91P_1_I92_1_T4), .i2(READ_ADD[5]), .i3(READ_ADD[4]), .o(N91P_1_I92_1_TC), .i0(READ_ADD[7]), .i1(READ_ADD[6]));
and2 N91P_1_I92_1_I34_1 (.o(N91P_1_I92_1_T5), .i0(READ_ADD[4]), .i1(N91P_1_I92_1_T4));
and2 N91P_1_I92_1_I32_1 (.o(N91P_1_UN_1_CB8CLE_I92_CEO), .i0(READ_ENABLE), .i1(N91P_1_I92_1_TC));
and2 N91P_1_I92_1_I30_1 (.o(N91P_1_I92_1_T2), .i0(READ_ADD[1]), .i1(READ_ADD[0]));
or2 N91P_1_I90_1_I23_1_I8_1_I5_1 (.o(N91P_1_I90_1_I23_1_MD[0]), .i0(N91P_1_I90_1_I23_1_I8_1_M1[0]), .i1(N91P_1_I90_1_I23_1_I8_1_M0[0]));
and2b1 N91P_1_I90_1_I23_1_I8_1_I7_1 (.o(N91P_1_I90_1_I23_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I90_1_I23_1_TQ[0]));
and2 N91P_1_I90_1_I23_1_I8_1_I6_1 (.o(N91P_1_I90_1_I23_1_I8_1_M1[0]), .i0(ADD_IN[17]), .i1(N91P_1_LD));
fdce N91P_1_I90_1_I23_1_I12_1 (.q(READ_ADD[17]), .d(N91P_1_I90_1_I23_1_MD[0]), .c(READ_CU), .ce(N91P_1_I90_1_I23_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I90_1_I23_1_I13_1 (.o(N91P_1_I90_1_I23_1_L_CE), .i0(N91P_1_UN_1_CB4CLE_I90_CE), .i1(N91P_1_LD));
xor2 N91P_1_I90_1_I23_1_I9_1 (.o(N91P_1_I90_1_I23_1_TQ[0]), .i0(READ_ADD[16]), .i1(READ_ADD[17]));
or2 N91P_1_I90_1_I22_1_I8_1_I5_1 (.o(N91P_1_I90_1_I22_1_MD[0]), .i0(N91P_1_I90_1_I22_1_I8_1_M1[0]), .i1(N91P_1_I90_1_I22_1_I8_1_M0[0]));
and2b1 N91P_1_I90_1_I22_1_I8_1_I7_1 (.o(N91P_1_I90_1_I22_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I90_1_I22_1_TQ[0]));
and2 N91P_1_I90_1_I22_1_I8_1_I6_1 (.o(N91P_1_I90_1_I22_1_I8_1_M1[0]), .i0(ADD_IN[16]), .i1(N91P_1_LD));
fdce N91P_1_I90_1_I22_1_I12_1 (.q(READ_ADD[16]), .d(N91P_1_I90_1_I22_1_MD[0]), .c(READ_CU), .ce(N91P_1_I90_1_I22_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I90_1_I22_1_I13_1 (.o(N91P_1_I90_1_I22_1_L_CE), .i0(N91P_1_UN_1_CB4CLE_I90_CE), .i1(N91P_1_LD));
xor2 N91P_1_I90_1_I22_1_I9_1 (.o(N91P_1_I90_1_I22_1_TQ[0]), .i0(XVDD), .i1(READ_ADD[16]));
or2 N91P_1_I90_1_I20_1_I8_1_I5_1 (.o(N91P_1_I90_1_I20_1_MD[0]), .i0(N91P_1_I90_1_I20_1_I8_1_M1[0]), .i1(N91P_1_I90_1_I20_1_I8_1_M0[0]));
and2b1 N91P_1_I90_1_I20_1_I8_1_I7_1 (.o(N91P_1_I90_1_I20_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I90_1_I20_1_TQ[0]));
and2 N91P_1_I90_1_I20_1_I8_1_I6_1 (.o(N91P_1_I90_1_I20_1_I8_1_M1[0]), .i0(ADD_IN[19]), .i1(N91P_1_LD));
fdce N91P_1_I90_1_I20_1_I12_1 (.q(READ_ADD[19]), .d(N91P_1_I90_1_I20_1_MD[0]), .c(READ_CU), .ce(N91P_1_I90_1_I20_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I90_1_I20_1_I13_1 (.o(N91P_1_I90_1_I20_1_L_CE), .i0(N91P_1_UN_1_CB4CLE_I90_CE), .i1(N91P_1_LD));
xor2 N91P_1_I90_1_I20_1_I9_1 (.o(N91P_1_I90_1_I20_1_TQ[0]), .i0(N91P_1_I90_1_T3), .i1(READ_ADD[19]));
or2 N91P_1_I90_1_I18_1_I8_1_I5_1 (.o(N91P_1_I90_1_I18_1_MD[0]), .i0(N91P_1_I90_1_I18_1_I8_1_M1[0]), .i1(N91P_1_I90_1_I18_1_I8_1_M0[0]));
and2b1 N91P_1_I90_1_I18_1_I8_1_I7_1 (.o(N91P_1_I90_1_I18_1_I8_1_M0[0]), .i0(N91P_1_LD), .i1(N91P_1_I90_1_I18_1_TQ[0]));
and2 N91P_1_I90_1_I18_1_I8_1_I6_1 (.o(N91P_1_I90_1_I18_1_I8_1_M1[0]), .i0(ADD_IN[18]), .i1(N91P_1_LD));
fdce N91P_1_I90_1_I18_1_I12_1 (.q(READ_ADD[18]), .d(N91P_1_I90_1_I18_1_MD[0]), .c(READ_CU), .ce(N91P_1_I90_1_I18_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N91P_1_I90_1_I18_1_I13_1 (.o(N91P_1_I90_1_I18_1_L_CE), .i0(N91P_1_UN_1_CB4CLE_I90_CE), .i1(N91P_1_LD));
xor2 N91P_1_I90_1_I18_1_I9_1 (.o(N91P_1_I90_1_I18_1_TQ[0]), .i0(N91P_1_I90_1_T2), .i1(READ_ADD[18]));
and3 N91P_1_I90_1_I21_1 (.i2(READ_ADD[16]), .o(N91P_1_I90_1_T3), .i0(READ_ADD[18]), .i1(READ_ADD[17]));
and4 N91P_1_I90_1_I19_1 (.i2(READ_ADD[18]), .i3(READ_ADD[19]), .o(N91P_1_I90_1_TC), .i0(READ_ADD[16]), .i1(READ_ADD[17]));
and2 N91P_1_I90_1_I24_1 (.o(N91P_1_I90_1_CEO), .i0(N91P_1_UN_1_CB4CLE_I90_CE), .i1(N91P_1_I90_1_TC));
and2 N91P_1_I90_1_I17_1 (.o(N91P_1_I90_1_T2), .i0(READ_ADD[17]), .i1(READ_ADD[16]));
buft N91P_1_I91_1_20 (.i(READ_ADD[19]), .o(XDT[19]), .t(REG_CNTROL[1]));
buft N91P_1_I91_1_19 (.t(REG_CNTROL[1]), .o(XDT[18]), .i(READ_ADD[18]));
buft N91P_1_I91_1_18 (.t(REG_CNTROL[1]), .o(XDT[17]), .i(READ_ADD[17]));
buft N91P_1_I91_1_17 (.t(REG_CNTROL[1]), .o(XDT[16]), .i(READ_ADD[16]));
buft N91P_1_I91_1_16 (.t(REG_CNTROL[1]), .o(XDT[15]), .i(READ_ADD[15]));
buft N91P_1_I91_1_15 (.t(REG_CNTROL[1]), .o(XDT[14]), .i(READ_ADD[14]));
buft N91P_1_I91_1_14 (.t(REG_CNTROL[1]), .o(XDT[13]), .i(READ_ADD[13]));
buft N91P_1_I91_1_13 (.t(REG_CNTROL[1]), .o(XDT[12]), .i(READ_ADD[12]));
buft N91P_1_I91_1_12 (.t(REG_CNTROL[1]), .o(XDT[11]), .i(READ_ADD[11]));
buft N91P_1_I91_1_11 (.t(REG_CNTROL[1]), .o(XDT[10]), .i(READ_ADD[10]));
buft N91P_1_I91_1_10 (.t(REG_CNTROL[1]), .o(XDT[9]), .i(READ_ADD[9]));
buft N91P_1_I91_1_9 (.t(REG_CNTROL[1]), .o(XDT[8]), .i(READ_ADD[8]));
buft N91P_1_I91_1_8 (.t(REG_CNTROL[1]), .o(XDT[7]), .i(READ_ADD[7]));
buft N91P_1_I91_1_7 (.t(REG_CNTROL[1]), .o(XDT[6]), .i(READ_ADD[6]));
buft N91P_1_I91_1_6 (.t(REG_CNTROL[1]), .o(XDT[5]), .i(READ_ADD[5]));
buft N91P_1_I91_1_5 (.t(REG_CNTROL[1]), .o(XDT[4]), .i(READ_ADD[4]));
buft N91P_1_I91_1_4 (.t(REG_CNTROL[1]), .o(XDT[3]), .i(READ_ADD[3]));
buft N91P_1_I91_1_3 (.t(REG_CNTROL[1]), .o(XDT[2]), .i(READ_ADD[2]));
buft N91P_1_I91_1_2 (.t(REG_CNTROL[1]), .o(XDT[1]), .i(READ_ADD[1]));
buft N91P_1_I91_1_1 (.t(REG_CNTROL[1]), .o(XDT[0]), .i(READ_ADD[0]));
inv N91P_1_94P_1 (.i(N_XREG_WR), .o(N91P_1_LD));
or2 N125P_1_I93_1_I44_1_I8_1_I5_1 (.o(N125P_1_I93_1_I44_1_MD[0]), .i0(N125P_1_I93_1_I44_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I44_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I44_1_I8_1_I7_1 (.o(N125P_1_I93_1_I44_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I44_1_TQ[0]));
and2 N125P_1_I93_1_I44_1_I8_1_I6_1 (.o(N125P_1_I93_1_I44_1_I8_1_M1[0]), .i0(ADD_IN[14]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I44_1_I12_1 (.q(WRITE_ADD[14]), .d(N125P_1_I93_1_I44_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I44_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I44_1_I13_1 (.o(N125P_1_I93_1_I44_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I44_1_I9_1 (.o(N125P_1_I93_1_I44_1_TQ[0]), .i0(N125P_1_I93_1_T6), .i1(WRITE_ADD[14]));
or2 N125P_1_I93_1_I43_1_I8_1_I5_1 (.o(N125P_1_I93_1_I43_1_MD[0]), .i0(N125P_1_I93_1_I43_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I43_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I43_1_I8_1_I7_1 (.o(N125P_1_I93_1_I43_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I43_1_TQ[0]));
and2 N125P_1_I93_1_I43_1_I8_1_I6_1 (.o(N125P_1_I93_1_I43_1_I8_1_M1[0]), .i0(ADD_IN[13]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I43_1_I12_1 (.q(WRITE_ADD[13]), .d(N125P_1_I93_1_I43_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I43_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I43_1_I13_1 (.o(N125P_1_I93_1_I43_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I43_1_I9_1 (.o(N125P_1_I93_1_I43_1_TQ[0]), .i0(N125P_1_I93_1_T5), .i1(WRITE_ADD[13]));
or2 N125P_1_I93_1_I39_1_I8_1_I5_1 (.o(N125P_1_I93_1_I39_1_MD[0]), .i0(N125P_1_I93_1_I39_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I39_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I39_1_I8_1_I7_1 (.o(N125P_1_I93_1_I39_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I39_1_TQ[0]));
and2 N125P_1_I93_1_I39_1_I8_1_I6_1 (.o(N125P_1_I93_1_I39_1_I8_1_M1[0]), .i0(ADD_IN[15]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I39_1_I12_1 (.q(WRITE_ADD[15]), .d(N125P_1_I93_1_I39_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I39_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I39_1_I13_1 (.o(N125P_1_I93_1_I39_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I39_1_I9_1 (.o(N125P_1_I93_1_I39_1_TQ[0]), .i0(N125P_1_I93_1_T7), .i1(WRITE_ADD[15]));
or2 N125P_1_I93_1_I36_1_I8_1_I5_1 (.o(N125P_1_I93_1_I36_1_MD[0]), .i0(N125P_1_I93_1_I36_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I36_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I36_1_I8_1_I7_1 (.o(N125P_1_I93_1_I36_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I36_1_TQ[0]));
and2 N125P_1_I93_1_I36_1_I8_1_I6_1 (.o(N125P_1_I93_1_I36_1_I8_1_M1[0]), .i0(ADD_IN[11]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I36_1_I12_1 (.q(WRITE_ADD[11]), .d(N125P_1_I93_1_I36_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I36_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I36_1_I13_1 (.o(N125P_1_I93_1_I36_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I36_1_I9_1 (.o(N125P_1_I93_1_I36_1_TQ[0]), .i0(N125P_1_I93_1_T3), .i1(WRITE_ADD[11]));
or2 N125P_1_I93_1_I35_1_I8_1_I5_1 (.o(N125P_1_I93_1_I35_1_MD[0]), .i0(N125P_1_I93_1_I35_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I35_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I35_1_I8_1_I7_1 (.o(N125P_1_I93_1_I35_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I35_1_TQ[0]));
and2 N125P_1_I93_1_I35_1_I8_1_I6_1 (.o(N125P_1_I93_1_I35_1_I8_1_M1[0]), .i0(ADD_IN[8]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I35_1_I12_1 (.q(WRITE_ADD[8]), .d(N125P_1_I93_1_I35_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I35_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I35_1_I13_1 (.o(N125P_1_I93_1_I35_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I35_1_I9_1 (.o(N125P_1_I93_1_I35_1_TQ[0]), .i0(XVDD), .i1(WRITE_ADD[8]));
or2 N125P_1_I93_1_I31_1_I8_1_I5_1 (.o(N125P_1_I93_1_I31_1_MD[0]), .i0(N125P_1_I93_1_I31_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I31_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I31_1_I8_1_I7_1 (.o(N125P_1_I93_1_I31_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I31_1_TQ[0]));
and2 N125P_1_I93_1_I31_1_I8_1_I6_1 (.o(N125P_1_I93_1_I31_1_I8_1_M1[0]), .i0(ADD_IN[9]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I31_1_I12_1 (.q(WRITE_ADD[9]), .d(N125P_1_I93_1_I31_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I31_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I31_1_I13_1 (.o(N125P_1_I93_1_I31_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I31_1_I9_1 (.o(N125P_1_I93_1_I31_1_TQ[0]), .i0(WRITE_ADD[8]), .i1(WRITE_ADD[9]));
or2 N125P_1_I93_1_I26_1_I8_1_I5_1 (.o(N125P_1_I93_1_I26_1_MD[0]), .i0(N125P_1_I93_1_I26_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I26_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I26_1_I8_1_I7_1 (.o(N125P_1_I93_1_I26_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I26_1_TQ[0]));
and2 N125P_1_I93_1_I26_1_I8_1_I6_1 (.o(N125P_1_I93_1_I26_1_I8_1_M1[0]), .i0(ADD_IN[10]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I26_1_I12_1 (.q(WRITE_ADD[10]), .d(N125P_1_I93_1_I26_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I26_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I26_1_I13_1 (.o(N125P_1_I93_1_I26_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I26_1_I9_1 (.o(N125P_1_I93_1_I26_1_TQ[0]), .i0(N125P_1_I93_1_T2), .i1(WRITE_ADD[10]));
or2 N125P_1_I93_1_I25_1_I8_1_I5_1 (.o(N125P_1_I93_1_I25_1_MD[0]), .i0(N125P_1_I93_1_I25_1_I8_1_M1[0]), .i1(N125P_1_I93_1_I25_1_I8_1_M0[0]));
and2b1 N125P_1_I93_1_I25_1_I8_1_I7_1 (.o(N125P_1_I93_1_I25_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I93_1_I25_1_TQ[0]));
and2 N125P_1_I93_1_I25_1_I8_1_I6_1 (.o(N125P_1_I93_1_I25_1_I8_1_M1[0]), .i0(ADD_IN[12]), .i1(N125P_1_LD));
fdce N125P_1_I93_1_I25_1_I12_1 (.q(WRITE_ADD[12]), .d(N125P_1_I93_1_I25_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I93_1_I25_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I93_1_I25_1_I13_1 (.o(N125P_1_I93_1_I25_1_L_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_LD));
xor2 N125P_1_I93_1_I25_1_I9_1 (.o(N125P_1_I93_1_I25_1_TQ[0]), .i0(N125P_1_I93_1_T4), .i1(WRITE_ADD[12]));
and3 N125P_1_I93_1_I29_1 (.i2(WRITE_ADD[8]), .o(N125P_1_I93_1_T3), .i0(WRITE_ADD[10]), .i1(WRITE_ADD[9]));
and3 N125P_1_I93_1_I27_1 (.i2(N125P_1_I93_1_T4), .o(N125P_1_I93_1_T6), .i0(WRITE_ADD[13]), .i1(WRITE_ADD[12]));
and4 N125P_1_I93_1_I38_1 (.i2(WRITE_ADD[9]), .i3(WRITE_ADD[8]), .o(N125P_1_I93_1_T4), .i0(WRITE_ADD[11]), .i1(WRITE_ADD[10]));
and4 N125P_1_I93_1_I33_1 (.i2(WRITE_ADD[12]), .i3(N125P_1_I93_1_T4), .o(N125P_1_I93_1_T7), .i0(WRITE_ADD[14]), .i1(WRITE_ADD[13]));
and5 N125P_1_I93_1_I37_1 (.i4(N125P_1_I93_1_T4), .i2(WRITE_ADD[13]), .i3(WRITE_ADD[12]), .o(N125P_1_I93_1_TC), .i0(WRITE_ADD[15]), .i1(WRITE_ADD[14]));
and2 N125P_1_I93_1_I34_1 (.o(N125P_1_I93_1_T5), .i0(WRITE_ADD[12]), .i1(N125P_1_I93_1_T4));
and2 N125P_1_I93_1_I32_1 (.o(N125P_1_UN_1_CB4CLE_I90_CE), .i0(N125P_1_UN_1_CB8CLE_I92_CEO), .i1(N125P_1_I93_1_TC));
and2 N125P_1_I93_1_I30_1 (.o(N125P_1_I93_1_T2), .i0(WRITE_ADD[9]), .i1(WRITE_ADD[8]));
or2 N125P_1_I92_1_I44_1_I8_1_I5_1 (.o(N125P_1_I92_1_I44_1_MD[0]), .i0(N125P_1_I92_1_I44_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I44_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I44_1_I8_1_I7_1 (.o(N125P_1_I92_1_I44_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I44_1_TQ[0]));
and2 N125P_1_I92_1_I44_1_I8_1_I6_1 (.o(N125P_1_I92_1_I44_1_I8_1_M1[0]), .i0(ADD_IN[6]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I44_1_I12_1 (.q(WRITE_ADD[6]), .d(N125P_1_I92_1_I44_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I44_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I44_1_I13_1 (.o(N125P_1_I92_1_I44_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I44_1_I9_1 (.o(N125P_1_I92_1_I44_1_TQ[0]), .i0(N125P_1_I92_1_T6), .i1(WRITE_ADD[6]));
or2 N125P_1_I92_1_I43_1_I8_1_I5_1 (.o(N125P_1_I92_1_I43_1_MD[0]), .i0(N125P_1_I92_1_I43_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I43_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I43_1_I8_1_I7_1 (.o(N125P_1_I92_1_I43_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I43_1_TQ[0]));
and2 N125P_1_I92_1_I43_1_I8_1_I6_1 (.o(N125P_1_I92_1_I43_1_I8_1_M1[0]), .i0(ADD_IN[5]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I43_1_I12_1 (.q(WRITE_ADD[5]), .d(N125P_1_I92_1_I43_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I43_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I43_1_I13_1 (.o(N125P_1_I92_1_I43_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I43_1_I9_1 (.o(N125P_1_I92_1_I43_1_TQ[0]), .i0(N125P_1_I92_1_T5), .i1(WRITE_ADD[5]));
or2 N125P_1_I92_1_I39_1_I8_1_I5_1 (.o(N125P_1_I92_1_I39_1_MD[0]), .i0(N125P_1_I92_1_I39_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I39_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I39_1_I8_1_I7_1 (.o(N125P_1_I92_1_I39_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I39_1_TQ[0]));
and2 N125P_1_I92_1_I39_1_I8_1_I6_1 (.o(N125P_1_I92_1_I39_1_I8_1_M1[0]), .i0(ADD_IN[7]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I39_1_I12_1 (.q(WRITE_ADD[7]), .d(N125P_1_I92_1_I39_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I39_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I39_1_I13_1 (.o(N125P_1_I92_1_I39_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I39_1_I9_1 (.o(N125P_1_I92_1_I39_1_TQ[0]), .i0(N125P_1_I92_1_T7), .i1(WRITE_ADD[7]));
or2 N125P_1_I92_1_I36_1_I8_1_I5_1 (.o(N125P_1_I92_1_I36_1_MD[0]), .i0(N125P_1_I92_1_I36_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I36_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I36_1_I8_1_I7_1 (.o(N125P_1_I92_1_I36_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I36_1_TQ[0]));
and2 N125P_1_I92_1_I36_1_I8_1_I6_1 (.o(N125P_1_I92_1_I36_1_I8_1_M1[0]), .i0(ADD_IN[3]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I36_1_I12_1 (.q(WRITE_ADD[3]), .d(N125P_1_I92_1_I36_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I36_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I36_1_I13_1 (.o(N125P_1_I92_1_I36_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I36_1_I9_1 (.o(N125P_1_I92_1_I36_1_TQ[0]), .i0(N125P_1_I92_1_T3), .i1(WRITE_ADD[3]));
or2 N125P_1_I92_1_I35_1_I8_1_I5_1 (.o(N125P_1_I92_1_I35_1_MD[0]), .i0(N125P_1_I92_1_I35_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I35_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I35_1_I8_1_I7_1 (.o(N125P_1_I92_1_I35_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I35_1_TQ[0]));
and2 N125P_1_I92_1_I35_1_I8_1_I6_1 (.o(N125P_1_I92_1_I35_1_I8_1_M1[0]), .i0(ADD_IN[0]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I35_1_I12_1 (.q(WRITE_ADD[0]), .d(N125P_1_I92_1_I35_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I35_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I35_1_I13_1 (.o(N125P_1_I92_1_I35_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I35_1_I9_1 (.o(N125P_1_I92_1_I35_1_TQ[0]), .i0(XVDD), .i1(WRITE_ADD[0]));
or2 N125P_1_I92_1_I31_1_I8_1_I5_1 (.o(N125P_1_I92_1_I31_1_MD[0]), .i0(N125P_1_I92_1_I31_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I31_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I31_1_I8_1_I7_1 (.o(N125P_1_I92_1_I31_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I31_1_TQ[0]));
and2 N125P_1_I92_1_I31_1_I8_1_I6_1 (.o(N125P_1_I92_1_I31_1_I8_1_M1[0]), .i0(ADD_IN[1]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I31_1_I12_1 (.q(WRITE_ADD[1]), .d(N125P_1_I92_1_I31_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I31_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I31_1_I13_1 (.o(N125P_1_I92_1_I31_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I31_1_I9_1 (.o(N125P_1_I92_1_I31_1_TQ[0]), .i0(WRITE_ADD[0]), .i1(WRITE_ADD[1]));
or2 N125P_1_I92_1_I26_1_I8_1_I5_1 (.o(N125P_1_I92_1_I26_1_MD[0]), .i0(N125P_1_I92_1_I26_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I26_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I26_1_I8_1_I7_1 (.o(N125P_1_I92_1_I26_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I26_1_TQ[0]));
and2 N125P_1_I92_1_I26_1_I8_1_I6_1 (.o(N125P_1_I92_1_I26_1_I8_1_M1[0]), .i0(ADD_IN[2]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I26_1_I12_1 (.q(WRITE_ADD[2]), .d(N125P_1_I92_1_I26_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I26_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I26_1_I13_1 (.o(N125P_1_I92_1_I26_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I26_1_I9_1 (.o(N125P_1_I92_1_I26_1_TQ[0]), .i0(N125P_1_I92_1_T2), .i1(WRITE_ADD[2]));
or2 N125P_1_I92_1_I25_1_I8_1_I5_1 (.o(N125P_1_I92_1_I25_1_MD[0]), .i0(N125P_1_I92_1_I25_1_I8_1_M1[0]), .i1(N125P_1_I92_1_I25_1_I8_1_M0[0]));
and2b1 N125P_1_I92_1_I25_1_I8_1_I7_1 (.o(N125P_1_I92_1_I25_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I92_1_I25_1_TQ[0]));
and2 N125P_1_I92_1_I25_1_I8_1_I6_1 (.o(N125P_1_I92_1_I25_1_I8_1_M1[0]), .i0(ADD_IN[4]), .i1(N125P_1_LD));
fdce N125P_1_I92_1_I25_1_I12_1 (.q(WRITE_ADD[4]), .d(N125P_1_I92_1_I25_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I92_1_I25_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I92_1_I25_1_I13_1 (.o(N125P_1_I92_1_I25_1_L_CE), .i0(WRITE_ENABLE), .i1(N125P_1_LD));
xor2 N125P_1_I92_1_I25_1_I9_1 (.o(N125P_1_I92_1_I25_1_TQ[0]), .i0(N125P_1_I92_1_T4), .i1(WRITE_ADD[4]));
and3 N125P_1_I92_1_I29_1 (.i2(WRITE_ADD[0]), .o(N125P_1_I92_1_T3), .i0(WRITE_ADD[2]), .i1(WRITE_ADD[1]));
and3 N125P_1_I92_1_I27_1 (.i2(N125P_1_I92_1_T4), .o(N125P_1_I92_1_T6), .i0(WRITE_ADD[5]), .i1(WRITE_ADD[4]));
and4 N125P_1_I92_1_I38_1 (.i2(WRITE_ADD[1]), .i3(WRITE_ADD[0]), .o(N125P_1_I92_1_T4), .i0(WRITE_ADD[3]), .i1(WRITE_ADD[2]));
and4 N125P_1_I92_1_I33_1 (.i2(WRITE_ADD[4]), .i3(N125P_1_I92_1_T4), .o(N125P_1_I92_1_T7), .i0(WRITE_ADD[6]), .i1(WRITE_ADD[5]));
and5 N125P_1_I92_1_I37_1 (.i4(N125P_1_I92_1_T4), .i2(WRITE_ADD[5]), .i3(WRITE_ADD[4]), .o(N125P_1_I92_1_TC), .i0(WRITE_ADD[7]), .i1(WRITE_ADD[6]));
and2 N125P_1_I92_1_I34_1 (.o(N125P_1_I92_1_T5), .i0(WRITE_ADD[4]), .i1(N125P_1_I92_1_T4));
and2 N125P_1_I92_1_I32_1 (.o(N125P_1_UN_1_CB8CLE_I92_CEO), .i0(WRITE_ENABLE), .i1(N125P_1_I92_1_TC));
and2 N125P_1_I92_1_I30_1 (.o(N125P_1_I92_1_T2), .i0(WRITE_ADD[1]), .i1(WRITE_ADD[0]));
or2 N125P_1_I90_1_I23_1_I8_1_I5_1 (.o(N125P_1_I90_1_I23_1_MD[0]), .i0(N125P_1_I90_1_I23_1_I8_1_M1[0]), .i1(N125P_1_I90_1_I23_1_I8_1_M0[0]));
and2b1 N125P_1_I90_1_I23_1_I8_1_I7_1 (.o(N125P_1_I90_1_I23_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I90_1_I23_1_TQ[0]));
and2 N125P_1_I90_1_I23_1_I8_1_I6_1 (.o(N125P_1_I90_1_I23_1_I8_1_M1[0]), .i0(ADD_IN[17]), .i1(N125P_1_LD));
fdce N125P_1_I90_1_I23_1_I12_1 (.q(WRITE_ADD[17]), .d(N125P_1_I90_1_I23_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I90_1_I23_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I90_1_I23_1_I13_1 (.o(N125P_1_I90_1_I23_1_L_CE), .i0(N125P_1_UN_1_CB4CLE_I90_CE), .i1(N125P_1_LD));
xor2 N125P_1_I90_1_I23_1_I9_1 (.o(N125P_1_I90_1_I23_1_TQ[0]), .i0(WRITE_ADD[16]), .i1(WRITE_ADD[17]));
or2 N125P_1_I90_1_I22_1_I8_1_I5_1 (.o(N125P_1_I90_1_I22_1_MD[0]), .i0(N125P_1_I90_1_I22_1_I8_1_M1[0]), .i1(N125P_1_I90_1_I22_1_I8_1_M0[0]));
and2b1 N125P_1_I90_1_I22_1_I8_1_I7_1 (.o(N125P_1_I90_1_I22_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I90_1_I22_1_TQ[0]));
and2 N125P_1_I90_1_I22_1_I8_1_I6_1 (.o(N125P_1_I90_1_I22_1_I8_1_M1[0]), .i0(ADD_IN[16]), .i1(N125P_1_LD));
fdce N125P_1_I90_1_I22_1_I12_1 (.q(WRITE_ADD[16]), .d(N125P_1_I90_1_I22_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I90_1_I22_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I90_1_I22_1_I13_1 (.o(N125P_1_I90_1_I22_1_L_CE), .i0(N125P_1_UN_1_CB4CLE_I90_CE), .i1(N125P_1_LD));
xor2 N125P_1_I90_1_I22_1_I9_1 (.o(N125P_1_I90_1_I22_1_TQ[0]), .i0(XVDD), .i1(WRITE_ADD[16]));
or2 N125P_1_I90_1_I20_1_I8_1_I5_1 (.o(N125P_1_I90_1_I20_1_MD[0]), .i0(N125P_1_I90_1_I20_1_I8_1_M1[0]), .i1(N125P_1_I90_1_I20_1_I8_1_M0[0]));
and2b1 N125P_1_I90_1_I20_1_I8_1_I7_1 (.o(N125P_1_I90_1_I20_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I90_1_I20_1_TQ[0]));
and2 N125P_1_I90_1_I20_1_I8_1_I6_1 (.o(N125P_1_I90_1_I20_1_I8_1_M1[0]), .i0(ADD_IN[19]), .i1(N125P_1_LD));
fdce N125P_1_I90_1_I20_1_I12_1 (.q(WRITE_ADD[19]), .d(N125P_1_I90_1_I20_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I90_1_I20_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I90_1_I20_1_I13_1 (.o(N125P_1_I90_1_I20_1_L_CE), .i0(N125P_1_UN_1_CB4CLE_I90_CE), .i1(N125P_1_LD));
xor2 N125P_1_I90_1_I20_1_I9_1 (.o(N125P_1_I90_1_I20_1_TQ[0]), .i0(N125P_1_I90_1_T3), .i1(WRITE_ADD[19]));
or2 N125P_1_I90_1_I18_1_I8_1_I5_1 (.o(N125P_1_I90_1_I18_1_MD[0]), .i0(N125P_1_I90_1_I18_1_I8_1_M1[0]), .i1(N125P_1_I90_1_I18_1_I8_1_M0[0]));
and2b1 N125P_1_I90_1_I18_1_I8_1_I7_1 (.o(N125P_1_I90_1_I18_1_I8_1_M0[0]), .i0(N125P_1_LD), .i1(N125P_1_I90_1_I18_1_TQ[0]));
and2 N125P_1_I90_1_I18_1_I8_1_I6_1 (.o(N125P_1_I90_1_I18_1_I8_1_M1[0]), .i0(ADD_IN[18]), .i1(N125P_1_LD));
fdce N125P_1_I90_1_I18_1_I12_1 (.q(WRITE_ADD[18]), .d(N125P_1_I90_1_I18_1_MD[0]), .c(WRITE_CU), .ce(N125P_1_I90_1_I18_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N125P_1_I90_1_I18_1_I13_1 (.o(N125P_1_I90_1_I18_1_L_CE), .i0(N125P_1_UN_1_CB4CLE_I90_CE), .i1(N125P_1_LD));
xor2 N125P_1_I90_1_I18_1_I9_1 (.o(N125P_1_I90_1_I18_1_TQ[0]), .i0(N125P_1_I90_1_T2), .i1(WRITE_ADD[18]));
and3 N125P_1_I90_1_I21_1 (.i2(WRITE_ADD[16]), .o(N125P_1_I90_1_T3), .i0(WRITE_ADD[18]), .i1(WRITE_ADD[17]));
and4 N125P_1_I90_1_I19_1 (.i2(WRITE_ADD[18]), .i3(WRITE_ADD[19]), .o(N125P_1_I90_1_TC), .i0(WRITE_ADD[16]), .i1(WRITE_ADD[17]));
and2 N125P_1_I90_1_I24_1 (.o(N125P_1_I90_1_CEO), .i0(N125P_1_UN_1_CB4CLE_I90_CE), .i1(N125P_1_I90_1_TC));
and2 N125P_1_I90_1_I17_1 (.o(N125P_1_I90_1_T2), .i0(WRITE_ADD[17]), .i1(WRITE_ADD[16]));
buft N125P_1_I91_1_20 (.i(WRITE_ADD[19]), .o(XDT[19]), .t(REG_CNTROL[0]));
buft N125P_1_I91_1_19 (.t(REG_CNTROL[0]), .o(XDT[18]), .i(WRITE_ADD[18]));
buft N125P_1_I91_1_18 (.t(REG_CNTROL[0]), .o(XDT[17]), .i(WRITE_ADD[17]));
buft N125P_1_I91_1_17 (.t(REG_CNTROL[0]), .o(XDT[16]), .i(WRITE_ADD[16]));
buft N125P_1_I91_1_16 (.t(REG_CNTROL[0]), .o(XDT[15]), .i(WRITE_ADD[15]));
buft N125P_1_I91_1_15 (.t(REG_CNTROL[0]), .o(XDT[14]), .i(WRITE_ADD[14]));
buft N125P_1_I91_1_14 (.t(REG_CNTROL[0]), .o(XDT[13]), .i(WRITE_ADD[13]));
buft N125P_1_I91_1_13 (.t(REG_CNTROL[0]), .o(XDT[12]), .i(WRITE_ADD[12]));
buft N125P_1_I91_1_12 (.t(REG_CNTROL[0]), .o(XDT[11]), .i(WRITE_ADD[11]));
buft N125P_1_I91_1_11 (.t(REG_CNTROL[0]), .o(XDT[10]), .i(WRITE_ADD[10]));
buft N125P_1_I91_1_10 (.t(REG_CNTROL[0]), .o(XDT[9]), .i(WRITE_ADD[9]));
buft N125P_1_I91_1_9 (.t(REG_CNTROL[0]), .o(XDT[8]), .i(WRITE_ADD[8]));
buft N125P_1_I91_1_8 (.t(REG_CNTROL[0]), .o(XDT[7]), .i(WRITE_ADD[7]));
buft N125P_1_I91_1_7 (.t(REG_CNTROL[0]), .o(XDT[6]), .i(WRITE_ADD[6]));
buft N125P_1_I91_1_6 (.t(REG_CNTROL[0]), .o(XDT[5]), .i(WRITE_ADD[5]));
buft N125P_1_I91_1_5 (.t(REG_CNTROL[0]), .o(XDT[4]), .i(WRITE_ADD[4]));
buft N125P_1_I91_1_4 (.t(REG_CNTROL[0]), .o(XDT[3]), .i(WRITE_ADD[3]));
buft N125P_1_I91_1_3 (.t(REG_CNTROL[0]), .o(XDT[2]), .i(WRITE_ADD[2]));
buft N125P_1_I91_1_2 (.t(REG_CNTROL[0]), .o(XDT[1]), .i(WRITE_ADD[1]));
buft N125P_1_I91_1_1 (.t(REG_CNTROL[0]), .o(XDT[0]), .i(WRITE_ADD[0]));
inv N125P_1_94P_1 (.i(N_XREG_WR), .o(N125P_1_LD));
or2 N107P_1_108P_1_I30_1_I6_1 (.o(N107P_1_108P_1_T1), .i0(N107P_1_108P_1_I30_1_M1[0]), .i1(N107P_1_108P_1_I30_1_M0[0]));
and2b2 N107P_1_108P_1_I30_1_I8_1 (.o(N107P_1_108P_1_I30_1_M0[0]), .i1(N_MEM_READ), .i0(N107P_1_POINTER_ADDRESS[0]));
and2 N107P_1_108P_1_I30_1_I5_1 (.o(N107P_1_108P_1_I30_1_M1[0]), .i0(N107P_1_POINTER_ADDRESS[0]), .i1(N_MEM_READ));
or2 N107P_1_108P_1_I49_1_I8_1_I5_1 (.o(N107P_1_108P_1_I49_1_MD[0]), .i0(N107P_1_108P_1_I49_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I49_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I49_1_I8_1_I7_1 (.o(N107P_1_108P_1_I49_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I49_1_TQ[0]));
and2 N107P_1_108P_1_I49_1_I8_1_I6_1 (.o(N107P_1_108P_1_I49_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[3]), .i1(XGND));
fdce N107P_1_108P_1_I49_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[3]), .d(N107P_1_108P_1_I49_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I49_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I49_1_I13_1 (.o(N107P_1_108P_1_I49_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I49_1_I9_1 (.o(N107P_1_108P_1_I49_1_TQ[0]), .i0(N107P_1_108P_1_T3), .i1(N107P_1_POINTER_ADDRESS[3]));
or2 N107P_1_108P_1_I46_1_I8_1_I5_1 (.o(N107P_1_108P_1_I46_1_MD[0]), .i0(N107P_1_108P_1_I46_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I46_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I46_1_I8_1_I7_1 (.o(N107P_1_108P_1_I46_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I46_1_TQ[0]));
and2 N107P_1_108P_1_I46_1_I8_1_I6_1 (.o(N107P_1_108P_1_I46_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[1]), .i1(XGND));
fdce N107P_1_108P_1_I46_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[1]), .d(N107P_1_108P_1_I46_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I46_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I46_1_I13_1 (.o(N107P_1_108P_1_I46_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I46_1_I9_1 (.o(N107P_1_108P_1_I46_1_TQ[0]), .i0(N107P_1_108P_1_T1), .i1(N107P_1_POINTER_ADDRESS[1]));
or2 N107P_1_108P_1_I42_1_I8_1_I5_1 (.o(N107P_1_108P_1_I42_1_MD[0]), .i0(N107P_1_108P_1_I42_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I42_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I42_1_I8_1_I7_1 (.o(N107P_1_108P_1_I42_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I42_1_TQ[0]));
and2 N107P_1_108P_1_I42_1_I8_1_I6_1 (.o(N107P_1_108P_1_I42_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[7]), .i1(XGND));
fdce N107P_1_108P_1_I42_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[7]), .d(N107P_1_108P_1_I42_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I42_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I42_1_I13_1 (.o(N107P_1_108P_1_I42_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I42_1_I9_1 (.o(N107P_1_108P_1_I42_1_TQ[0]), .i0(N107P_1_108P_1_T7), .i1(N107P_1_POINTER_ADDRESS[7]));
or2 N107P_1_108P_1_I43_1_I8_1_I5_1 (.o(N107P_1_108P_1_I43_1_MD[0]), .i0(N107P_1_108P_1_I43_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I43_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I43_1_I8_1_I7_1 (.o(N107P_1_108P_1_I43_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I43_1_TQ[0]));
and2 N107P_1_108P_1_I43_1_I8_1_I6_1 (.o(N107P_1_108P_1_I43_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[6]), .i1(XGND));
fdce N107P_1_108P_1_I43_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[6]), .d(N107P_1_108P_1_I43_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I43_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I43_1_I13_1 (.o(N107P_1_108P_1_I43_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I43_1_I9_1 (.o(N107P_1_108P_1_I43_1_TQ[0]), .i0(N107P_1_108P_1_T6), .i1(N107P_1_POINTER_ADDRESS[6]));
or2 N107P_1_108P_1_I35_1_I8_1_I5_1 (.o(N107P_1_108P_1_I35_1_MD[0]), .i0(N107P_1_108P_1_I35_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I35_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I35_1_I8_1_I7_1 (.o(N107P_1_108P_1_I35_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I35_1_TQ[0]));
and2 N107P_1_108P_1_I35_1_I8_1_I6_1 (.o(N107P_1_108P_1_I35_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[2]), .i1(XGND));
fdce N107P_1_108P_1_I35_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[2]), .d(N107P_1_108P_1_I35_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I35_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I35_1_I13_1 (.o(N107P_1_108P_1_I35_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I35_1_I9_1 (.o(N107P_1_108P_1_I35_1_TQ[0]), .i0(N107P_1_108P_1_T2), .i1(N107P_1_POINTER_ADDRESS[2]));
or2 N107P_1_108P_1_I34_1_I8_1_I5_1 (.o(N107P_1_108P_1_I34_1_MD[0]), .i0(N107P_1_108P_1_I34_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I34_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I34_1_I8_1_I7_1 (.o(N107P_1_108P_1_I34_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I34_1_TQ[0]));
and2 N107P_1_108P_1_I34_1_I8_1_I6_1 (.o(N107P_1_108P_1_I34_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[4]), .i1(XGND));
fdce N107P_1_108P_1_I34_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[4]), .d(N107P_1_108P_1_I34_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I34_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I34_1_I13_1 (.o(N107P_1_108P_1_I34_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I34_1_I9_1 (.o(N107P_1_108P_1_I34_1_TQ[0]), .i0(N107P_1_108P_1_T4), .i1(N107P_1_POINTER_ADDRESS[4]));
or2 N107P_1_108P_1_I31_1_I8_1_I5_1 (.o(N107P_1_108P_1_I31_1_MD[0]), .i0(N107P_1_108P_1_I31_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I31_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I31_1_I8_1_I7_1 (.o(N107P_1_108P_1_I31_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I31_1_TQ[0]));
and2 N107P_1_108P_1_I31_1_I8_1_I6_1 (.o(N107P_1_108P_1_I31_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[5]), .i1(XGND));
fdce N107P_1_108P_1_I31_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[5]), .d(N107P_1_108P_1_I31_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I31_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I31_1_I13_1 (.o(N107P_1_108P_1_I31_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I31_1_I9_1 (.o(N107P_1_108P_1_I31_1_TQ[0]), .i0(N107P_1_108P_1_T5), .i1(N107P_1_POINTER_ADDRESS[5]));
or2 N107P_1_108P_1_I29_1_I8_1_I5_1 (.o(N107P_1_108P_1_I29_1_MD[0]), .i0(N107P_1_108P_1_I29_1_I8_1_M1[0]), .i1(N107P_1_108P_1_I29_1_I8_1_M0[0]));
and2b1 N107P_1_108P_1_I29_1_I8_1_I7_1 (.o(N107P_1_108P_1_I29_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_108P_1_I29_1_TQ[0]));
and2 N107P_1_108P_1_I29_1_I8_1_I6_1 (.o(N107P_1_108P_1_I29_1_I8_1_M1[0]), .i0(N107P_1_108P_1_D[0]), .i1(XGND));
fdce N107P_1_108P_1_I29_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[0]), .d(N107P_1_108P_1_I29_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_108P_1_I29_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_108P_1_I29_1_I13_1 (.o(N107P_1_108P_1_I29_1_L_CE), .i0(XVDD), .i1(XGND));
xor2 N107P_1_108P_1_I29_1_I9_1 (.o(N107P_1_108P_1_I29_1_TQ[0]), .i0(XVDD), .i1(N107P_1_POINTER_ADDRESS[0]));
or2 N107P_1_108P_1_I57_1_I5_1 (.o(N107P_1_108P_1_TC), .i0(N107P_1_108P_1_I57_1_M1[0]), .i1(N107P_1_108P_1_I57_1_M0[0]));
and2b1 N107P_1_108P_1_I57_1_I7_1 (.o(N107P_1_108P_1_I57_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_108P_1_TC_DN));
and2 N107P_1_108P_1_I57_1_I6_1 (.o(N107P_1_108P_1_I57_1_M1[0]), .i0(N107P_1_108P_1_TC_UP), .i1(N_MEM_READ));
or2 N107P_1_108P_1_I56_1_I5_1 (.o(N107P_1_108P_1_T6), .i0(N107P_1_108P_1_I56_1_M1[0]), .i1(N107P_1_108P_1_I56_1_M0[0]));
and2b1 N107P_1_108P_1_I56_1_I7_1 (.o(N107P_1_108P_1_I56_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_108P_1_T6_DN));
and2 N107P_1_108P_1_I56_1_I6_1 (.o(N107P_1_108P_1_I56_1_M1[0]), .i0(N107P_1_108P_1_T6_UP), .i1(N_MEM_READ));
or2 N107P_1_108P_1_I41_1_I5_1 (.o(N107P_1_108P_1_T4), .i0(N107P_1_108P_1_I41_1_M1[0]), .i1(N107P_1_108P_1_I41_1_M0[0]));
and2b1 N107P_1_108P_1_I41_1_I7_1 (.o(N107P_1_108P_1_I41_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_108P_1_T4_DN));
and2 N107P_1_108P_1_I41_1_I6_1 (.o(N107P_1_108P_1_I41_1_M1[0]), .i0(N107P_1_108P_1_T4_UP), .i1(N_MEM_READ));
or2 N107P_1_108P_1_I40_1_I5_1 (.o(N107P_1_108P_1_T5), .i0(N107P_1_108P_1_I40_1_M1[0]), .i1(N107P_1_108P_1_I40_1_M0[0]));
and2b1 N107P_1_108P_1_I40_1_I7_1 (.o(N107P_1_108P_1_I40_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_108P_1_T5_DN));
and2 N107P_1_108P_1_I40_1_I6_1 (.o(N107P_1_108P_1_I40_1_M1[0]), .i0(N107P_1_108P_1_T5_UP), .i1(N_MEM_READ));
or2 N107P_1_108P_1_I44_1_I5_1 (.o(N107P_1_108P_1_T2), .i0(N107P_1_108P_1_I44_1_M1[0]), .i1(N107P_1_108P_1_I44_1_M0[0]));
and2b1 N107P_1_108P_1_I44_1_I7_1 (.o(N107P_1_108P_1_I44_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_108P_1_T2_DN));
and2 N107P_1_108P_1_I44_1_I6_1 (.o(N107P_1_108P_1_I44_1_M1[0]), .i0(N107P_1_108P_1_T2_UP), .i1(N_MEM_READ));
or2 N107P_1_108P_1_I36_1_I5_1 (.o(N107P_1_108P_1_T3), .i0(N107P_1_108P_1_I36_1_M1[0]), .i1(N107P_1_108P_1_I36_1_M0[0]));
and2b1 N107P_1_108P_1_I36_1_I7_1 (.o(N107P_1_108P_1_I36_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_108P_1_T3_DN));
and2 N107P_1_108P_1_I36_1_I6_1 (.o(N107P_1_108P_1_I36_1_M1[0]), .i0(N107P_1_108P_1_T3_UP), .i1(N_MEM_READ));
or2 N107P_1_108P_1_I27_1_I5_1 (.o(N107P_1_108P_1_T7), .i0(N107P_1_108P_1_I27_1_M1[0]), .i1(N107P_1_108P_1_I27_1_M0[0]));
and2b1 N107P_1_108P_1_I27_1_I7_1 (.o(N107P_1_108P_1_I27_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_108P_1_T7_DN));
and2 N107P_1_108P_1_I27_1_I6_1 (.o(N107P_1_108P_1_I27_1_M1[0]), .i0(N107P_1_108P_1_T7_UP), .i1(N_MEM_READ));
and3b2 N107P_1_108P_1_I53_1 (.i2(N107P_1_108P_1_T6), .o(N107P_1_108P_1_TC_DN), .i1(N107P_1_POINTER_ADDRESS[7]), .i0(N107P_1_POINTER_ADDRESS[6]));
and3b2 N107P_1_108P_1_I51_1 (.i2(N107P_1_108P_1_T3), .o(N107P_1_108P_1_T5_DN), .i1(N107P_1_POINTER_ADDRESS[4]), .i0(N107P_1_POINTER_ADDRESS[3]));
and4b3 N107P_1_108P_1_I26_1 (.i2(N107P_1_POINTER_ADDRESS[3]), .i3(N107P_1_108P_1_T3), .o(N107P_1_108P_1_T6_DN), .i1(N107P_1_POINTER_ADDRESS[5]), .i0(N107P_1_POINTER_ADDRESS[4]));
and3b3 N107P_1_108P_1_I45_1 (.i2(N107P_1_POINTER_ADDRESS[0]), .o(N107P_1_108P_1_T3_DN), .i1(N107P_1_POINTER_ADDRESS[2]), .i0(N107P_1_POINTER_ADDRESS[1]));
and2b2 N107P_1_108P_1_I37_1 (.o(N107P_1_108P_1_T2_DN), .i1(N107P_1_POINTER_ADDRESS[1]), .i0(N107P_1_POINTER_ADDRESS[0]));
and3 N107P_1_108P_1_I58_1 (.i2(N107P_1_POINTER_ADDRESS[0]), .o(N107P_1_108P_1_T3_UP), .i0(N107P_1_POINTER_ADDRESS[2]), .i1(N107P_1_POINTER_ADDRESS[1]));
and3 N107P_1_108P_1_I55_1 (.i2(N107P_1_108P_1_T3), .o(N107P_1_108P_1_T5_UP), .i0(N107P_1_POINTER_ADDRESS[4]), .i1(N107P_1_POINTER_ADDRESS[3]));
and3 N107P_1_108P_1_I47_1 (.i2(N107P_1_108P_1_T6), .o(N107P_1_108P_1_TC_UP), .i0(N107P_1_POINTER_ADDRESS[7]), .i1(N107P_1_POINTER_ADDRESS[6]));
and4 N107P_1_108P_1_I59_1 (.i2(N107P_1_POINTER_ADDRESS[3]), .i3(N107P_1_108P_1_T3), .o(N107P_1_108P_1_T6_UP), .i0(N107P_1_POINTER_ADDRESS[5]), .i1(N107P_1_POINTER_ADDRESS[4]));
and2b1 N107P_1_108P_1_I48_1 (.o(N107P_1_108P_1_T7_DN), .i0(N107P_1_POINTER_ADDRESS[6]), .i1(N107P_1_108P_1_T6));
and2b1 N107P_1_108P_1_I32_1 (.o(N107P_1_108P_1_T4_DN), .i0(N107P_1_POINTER_ADDRESS[3]), .i1(N107P_1_108P_1_T3));
and2 N107P_1_108P_1_I60_1 (.o(N107P_1_108P_1_T2_UP), .i0(N107P_1_POINTER_ADDRESS[1]), .i1(N107P_1_POINTER_ADDRESS[0]));
and2 N107P_1_108P_1_I54_1 (.o(N107P_1_UN_1_CB8CLED_107P_CE), .i0(XVDD), .i1(N107P_1_108P_1_TC));
and2 N107P_1_108P_1_I38_1 (.o(N107P_1_108P_1_T4_UP), .i0(N107P_1_POINTER_ADDRESS[3]), .i1(N107P_1_108P_1_T3));
and2 N107P_1_108P_1_I28_1 (.o(N107P_1_108P_1_T7_UP), .i0(N107P_1_POINTER_ADDRESS[6]), .i1(N107P_1_108P_1_T6));
or2 N107P_1_107P_1_I30_1_I6_1 (.o(N107P_1_107P_1_T1), .i0(N107P_1_107P_1_I30_1_M1[0]), .i1(N107P_1_107P_1_I30_1_M0[0]));
and2b2 N107P_1_107P_1_I30_1_I8_1 (.o(N107P_1_107P_1_I30_1_M0[0]), .i1(N_MEM_READ), .i0(N107P_1_POINTER_ADDRESS[8]));
and2 N107P_1_107P_1_I30_1_I5_1 (.o(N107P_1_107P_1_I30_1_M1[0]), .i0(N107P_1_POINTER_ADDRESS[8]), .i1(N_MEM_READ));
or2 N107P_1_107P_1_I49_1_I8_1_I5_1 (.o(N107P_1_107P_1_I49_1_MD[0]), .i0(N107P_1_107P_1_I49_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I49_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I49_1_I8_1_I7_1 (.o(N107P_1_107P_1_I49_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I49_1_TQ[0]));
and2 N107P_1_107P_1_I49_1_I8_1_I6_1 (.o(N107P_1_107P_1_I49_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[3]), .i1(XGND));
fdce N107P_1_107P_1_I49_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[11]), .d(N107P_1_107P_1_I49_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I49_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I49_1_I13_1 (.o(N107P_1_107P_1_I49_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I49_1_I9_1 (.o(N107P_1_107P_1_I49_1_TQ[0]), .i0(N107P_1_107P_1_T3), .i1(N107P_1_POINTER_ADDRESS[11]));
or2 N107P_1_107P_1_I46_1_I8_1_I5_1 (.o(N107P_1_107P_1_I46_1_MD[0]), .i0(N107P_1_107P_1_I46_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I46_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I46_1_I8_1_I7_1 (.o(N107P_1_107P_1_I46_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I46_1_TQ[0]));
and2 N107P_1_107P_1_I46_1_I8_1_I6_1 (.o(N107P_1_107P_1_I46_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[1]), .i1(XGND));
fdce N107P_1_107P_1_I46_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[9]), .d(N107P_1_107P_1_I46_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I46_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I46_1_I13_1 (.o(N107P_1_107P_1_I46_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I46_1_I9_1 (.o(N107P_1_107P_1_I46_1_TQ[0]), .i0(N107P_1_107P_1_T1), .i1(N107P_1_POINTER_ADDRESS[9]));
or2 N107P_1_107P_1_I42_1_I8_1_I5_1 (.o(N107P_1_107P_1_I42_1_MD[0]), .i0(N107P_1_107P_1_I42_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I42_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I42_1_I8_1_I7_1 (.o(N107P_1_107P_1_I42_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I42_1_TQ[0]));
and2 N107P_1_107P_1_I42_1_I8_1_I6_1 (.o(N107P_1_107P_1_I42_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[7]), .i1(XGND));
fdce N107P_1_107P_1_I42_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[15]), .d(N107P_1_107P_1_I42_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I42_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I42_1_I13_1 (.o(N107P_1_107P_1_I42_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I42_1_I9_1 (.o(N107P_1_107P_1_I42_1_TQ[0]), .i0(N107P_1_107P_1_T7), .i1(N107P_1_POINTER_ADDRESS[15]));
or2 N107P_1_107P_1_I43_1_I8_1_I5_1 (.o(N107P_1_107P_1_I43_1_MD[0]), .i0(N107P_1_107P_1_I43_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I43_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I43_1_I8_1_I7_1 (.o(N107P_1_107P_1_I43_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I43_1_TQ[0]));
and2 N107P_1_107P_1_I43_1_I8_1_I6_1 (.o(N107P_1_107P_1_I43_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[6]), .i1(XGND));
fdce N107P_1_107P_1_I43_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[14]), .d(N107P_1_107P_1_I43_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I43_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I43_1_I13_1 (.o(N107P_1_107P_1_I43_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I43_1_I9_1 (.o(N107P_1_107P_1_I43_1_TQ[0]), .i0(N107P_1_107P_1_T6), .i1(N107P_1_POINTER_ADDRESS[14]));
or2 N107P_1_107P_1_I35_1_I8_1_I5_1 (.o(N107P_1_107P_1_I35_1_MD[0]), .i0(N107P_1_107P_1_I35_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I35_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I35_1_I8_1_I7_1 (.o(N107P_1_107P_1_I35_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I35_1_TQ[0]));
and2 N107P_1_107P_1_I35_1_I8_1_I6_1 (.o(N107P_1_107P_1_I35_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[2]), .i1(XGND));
fdce N107P_1_107P_1_I35_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[10]), .d(N107P_1_107P_1_I35_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I35_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I35_1_I13_1 (.o(N107P_1_107P_1_I35_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I35_1_I9_1 (.o(N107P_1_107P_1_I35_1_TQ[0]), .i0(N107P_1_107P_1_T2), .i1(N107P_1_POINTER_ADDRESS[10]));
or2 N107P_1_107P_1_I34_1_I8_1_I5_1 (.o(N107P_1_107P_1_I34_1_MD[0]), .i0(N107P_1_107P_1_I34_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I34_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I34_1_I8_1_I7_1 (.o(N107P_1_107P_1_I34_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I34_1_TQ[0]));
and2 N107P_1_107P_1_I34_1_I8_1_I6_1 (.o(N107P_1_107P_1_I34_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[4]), .i1(XGND));
fdce N107P_1_107P_1_I34_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[12]), .d(N107P_1_107P_1_I34_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I34_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I34_1_I13_1 (.o(N107P_1_107P_1_I34_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I34_1_I9_1 (.o(N107P_1_107P_1_I34_1_TQ[0]), .i0(N107P_1_107P_1_T4), .i1(N107P_1_POINTER_ADDRESS[12]));
or2 N107P_1_107P_1_I31_1_I8_1_I5_1 (.o(N107P_1_107P_1_I31_1_MD[0]), .i0(N107P_1_107P_1_I31_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I31_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I31_1_I8_1_I7_1 (.o(N107P_1_107P_1_I31_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I31_1_TQ[0]));
and2 N107P_1_107P_1_I31_1_I8_1_I6_1 (.o(N107P_1_107P_1_I31_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[5]), .i1(XGND));
fdce N107P_1_107P_1_I31_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[13]), .d(N107P_1_107P_1_I31_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I31_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I31_1_I13_1 (.o(N107P_1_107P_1_I31_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I31_1_I9_1 (.o(N107P_1_107P_1_I31_1_TQ[0]), .i0(N107P_1_107P_1_T5), .i1(N107P_1_POINTER_ADDRESS[13]));
or2 N107P_1_107P_1_I29_1_I8_1_I5_1 (.o(N107P_1_107P_1_I29_1_MD[0]), .i0(N107P_1_107P_1_I29_1_I8_1_M1[0]), .i1(N107P_1_107P_1_I29_1_I8_1_M0[0]));
and2b1 N107P_1_107P_1_I29_1_I8_1_I7_1 (.o(N107P_1_107P_1_I29_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_107P_1_I29_1_TQ[0]));
and2 N107P_1_107P_1_I29_1_I8_1_I6_1 (.o(N107P_1_107P_1_I29_1_I8_1_M1[0]), .i0(N107P_1_107P_1_D[0]), .i1(XGND));
fdce N107P_1_107P_1_I29_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[8]), .d(N107P_1_107P_1_I29_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_107P_1_I29_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_107P_1_I29_1_I13_1 (.o(N107P_1_107P_1_I29_1_L_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(XGND));
xor2 N107P_1_107P_1_I29_1_I9_1 (.o(N107P_1_107P_1_I29_1_TQ[0]), .i0(XVDD), .i1(N107P_1_POINTER_ADDRESS[8]));
or2 N107P_1_107P_1_I57_1_I5_1 (.o(N107P_1_107P_1_TC), .i0(N107P_1_107P_1_I57_1_M1[0]), .i1(N107P_1_107P_1_I57_1_M0[0]));
and2b1 N107P_1_107P_1_I57_1_I7_1 (.o(N107P_1_107P_1_I57_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_107P_1_TC_DN));
and2 N107P_1_107P_1_I57_1_I6_1 (.o(N107P_1_107P_1_I57_1_M1[0]), .i0(N107P_1_107P_1_TC_UP), .i1(N_MEM_READ));
or2 N107P_1_107P_1_I56_1_I5_1 (.o(N107P_1_107P_1_T6), .i0(N107P_1_107P_1_I56_1_M1[0]), .i1(N107P_1_107P_1_I56_1_M0[0]));
and2b1 N107P_1_107P_1_I56_1_I7_1 (.o(N107P_1_107P_1_I56_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_107P_1_T6_DN));
and2 N107P_1_107P_1_I56_1_I6_1 (.o(N107P_1_107P_1_I56_1_M1[0]), .i0(N107P_1_107P_1_T6_UP), .i1(N_MEM_READ));
or2 N107P_1_107P_1_I41_1_I5_1 (.o(N107P_1_107P_1_T4), .i0(N107P_1_107P_1_I41_1_M1[0]), .i1(N107P_1_107P_1_I41_1_M0[0]));
and2b1 N107P_1_107P_1_I41_1_I7_1 (.o(N107P_1_107P_1_I41_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_107P_1_T4_DN));
and2 N107P_1_107P_1_I41_1_I6_1 (.o(N107P_1_107P_1_I41_1_M1[0]), .i0(N107P_1_107P_1_T4_UP), .i1(N_MEM_READ));
or2 N107P_1_107P_1_I40_1_I5_1 (.o(N107P_1_107P_1_T5), .i0(N107P_1_107P_1_I40_1_M1[0]), .i1(N107P_1_107P_1_I40_1_M0[0]));
and2b1 N107P_1_107P_1_I40_1_I7_1 (.o(N107P_1_107P_1_I40_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_107P_1_T5_DN));
and2 N107P_1_107P_1_I40_1_I6_1 (.o(N107P_1_107P_1_I40_1_M1[0]), .i0(N107P_1_107P_1_T5_UP), .i1(N_MEM_READ));
or2 N107P_1_107P_1_I44_1_I5_1 (.o(N107P_1_107P_1_T2), .i0(N107P_1_107P_1_I44_1_M1[0]), .i1(N107P_1_107P_1_I44_1_M0[0]));
and2b1 N107P_1_107P_1_I44_1_I7_1 (.o(N107P_1_107P_1_I44_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_107P_1_T2_DN));
and2 N107P_1_107P_1_I44_1_I6_1 (.o(N107P_1_107P_1_I44_1_M1[0]), .i0(N107P_1_107P_1_T2_UP), .i1(N_MEM_READ));
or2 N107P_1_107P_1_I36_1_I5_1 (.o(N107P_1_107P_1_T3), .i0(N107P_1_107P_1_I36_1_M1[0]), .i1(N107P_1_107P_1_I36_1_M0[0]));
and2b1 N107P_1_107P_1_I36_1_I7_1 (.o(N107P_1_107P_1_I36_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_107P_1_T3_DN));
and2 N107P_1_107P_1_I36_1_I6_1 (.o(N107P_1_107P_1_I36_1_M1[0]), .i0(N107P_1_107P_1_T3_UP), .i1(N_MEM_READ));
or2 N107P_1_107P_1_I27_1_I5_1 (.o(N107P_1_107P_1_T7), .i0(N107P_1_107P_1_I27_1_M1[0]), .i1(N107P_1_107P_1_I27_1_M0[0]));
and2b1 N107P_1_107P_1_I27_1_I7_1 (.o(N107P_1_107P_1_I27_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_107P_1_T7_DN));
and2 N107P_1_107P_1_I27_1_I6_1 (.o(N107P_1_107P_1_I27_1_M1[0]), .i0(N107P_1_107P_1_T7_UP), .i1(N_MEM_READ));
and3b2 N107P_1_107P_1_I53_1 (.i2(N107P_1_107P_1_T6), .o(N107P_1_107P_1_TC_DN), .i1(N107P_1_POINTER_ADDRESS[15]), .i0(N107P_1_POINTER_ADDRESS[14]));
and3b2 N107P_1_107P_1_I51_1 (.i2(N107P_1_107P_1_T3), .o(N107P_1_107P_1_T5_DN), .i1(N107P_1_POINTER_ADDRESS[12]), .i0(N107P_1_POINTER_ADDRESS[11]));
and4b3 N107P_1_107P_1_I26_1 (.i2(N107P_1_POINTER_ADDRESS[11]), .i3(N107P_1_107P_1_T3), .o(N107P_1_107P_1_T6_DN), .i1(N107P_1_POINTER_ADDRESS[13]), .i0(N107P_1_POINTER_ADDRESS[12]));
and3b3 N107P_1_107P_1_I45_1 (.i2(N107P_1_POINTER_ADDRESS[8]), .o(N107P_1_107P_1_T3_DN), .i1(N107P_1_POINTER_ADDRESS[10]), .i0(N107P_1_POINTER_ADDRESS[9]));
and2b2 N107P_1_107P_1_I37_1 (.o(N107P_1_107P_1_T2_DN), .i1(N107P_1_POINTER_ADDRESS[9]), .i0(N107P_1_POINTER_ADDRESS[8]));
and3 N107P_1_107P_1_I58_1 (.i2(N107P_1_POINTER_ADDRESS[8]), .o(N107P_1_107P_1_T3_UP), .i0(N107P_1_POINTER_ADDRESS[10]), .i1(N107P_1_POINTER_ADDRESS[9]));
and3 N107P_1_107P_1_I55_1 (.i2(N107P_1_107P_1_T3), .o(N107P_1_107P_1_T5_UP), .i0(N107P_1_POINTER_ADDRESS[12]), .i1(N107P_1_POINTER_ADDRESS[11]));
and3 N107P_1_107P_1_I47_1 (.i2(N107P_1_107P_1_T6), .o(N107P_1_107P_1_TC_UP), .i0(N107P_1_POINTER_ADDRESS[15]), .i1(N107P_1_POINTER_ADDRESS[14]));
and4 N107P_1_107P_1_I59_1 (.i2(N107P_1_POINTER_ADDRESS[11]), .i3(N107P_1_107P_1_T3), .o(N107P_1_107P_1_T6_UP), .i0(N107P_1_POINTER_ADDRESS[13]), .i1(N107P_1_POINTER_ADDRESS[12]));
and2b1 N107P_1_107P_1_I48_1 (.o(N107P_1_107P_1_T7_DN), .i0(N107P_1_POINTER_ADDRESS[14]), .i1(N107P_1_107P_1_T6));
and2b1 N107P_1_107P_1_I32_1 (.o(N107P_1_107P_1_T4_DN), .i0(N107P_1_POINTER_ADDRESS[11]), .i1(N107P_1_107P_1_T3));
and2 N107P_1_107P_1_I60_1 (.o(N107P_1_107P_1_T2_UP), .i0(N107P_1_POINTER_ADDRESS[9]), .i1(N107P_1_POINTER_ADDRESS[8]));
and2 N107P_1_107P_1_I54_1 (.o(N107P_1_UN_1_CB4CLED_100P_CE), .i0(N107P_1_UN_1_CB8CLED_107P_CE), .i1(N107P_1_107P_1_TC));
and2 N107P_1_107P_1_I38_1 (.o(N107P_1_107P_1_T4_UP), .i0(N107P_1_POINTER_ADDRESS[11]), .i1(N107P_1_107P_1_T3));
and2 N107P_1_107P_1_I28_1 (.o(N107P_1_107P_1_T7_UP), .i0(N107P_1_POINTER_ADDRESS[14]), .i1(N107P_1_107P_1_T6));
or2 N107P_1_100P_1_I27_1_I6_1 (.o(N107P_1_100P_1_T1), .i0(N107P_1_100P_1_I27_1_M1[0]), .i1(N107P_1_100P_1_I27_1_M0[0]));
and2b2 N107P_1_100P_1_I27_1_I8_1 (.o(N107P_1_100P_1_I27_1_M0[0]), .i1(N_MEM_READ), .i0(N107P_1_POINTER_ADDRESS[16]));
and2 N107P_1_100P_1_I27_1_I5_1 (.o(N107P_1_100P_1_I27_1_M1[0]), .i0(N107P_1_POINTER_ADDRESS[16]), .i1(N_MEM_READ));
or2 N107P_1_100P_1_I26_1_I8_1_I5_1 (.o(N107P_1_100P_1_I26_1_MD[0]), .i0(N107P_1_100P_1_I26_1_I8_1_M1[0]), .i1(N107P_1_100P_1_I26_1_I8_1_M0[0]));
and2b1 N107P_1_100P_1_I26_1_I8_1_I7_1 (.o(N107P_1_100P_1_I26_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_100P_1_I26_1_TQ[0]));
and2 N107P_1_100P_1_I26_1_I8_1_I6_1 (.o(N107P_1_100P_1_I26_1_I8_1_M1[0]), .i0(N107P_1_100P_1_D1), .i1(XGND));
fdce N107P_1_100P_1_I26_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[17]), .d(N107P_1_100P_1_I26_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_100P_1_I26_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_100P_1_I26_1_I13_1 (.o(N107P_1_100P_1_I26_1_L_CE), .i0(N107P_1_UN_1_CB4CLED_100P_CE), .i1(XGND));
xor2 N107P_1_100P_1_I26_1_I9_1 (.o(N107P_1_100P_1_I26_1_TQ[0]), .i0(N107P_1_100P_1_T1), .i1(N107P_1_POINTER_ADDRESS[17]));
or2 N107P_1_100P_1_I25_1_I8_1_I5_1 (.o(N107P_1_100P_1_I25_1_MD[0]), .i0(N107P_1_100P_1_I25_1_I8_1_M1[0]), .i1(N107P_1_100P_1_I25_1_I8_1_M0[0]));
and2b1 N107P_1_100P_1_I25_1_I8_1_I7_1 (.o(N107P_1_100P_1_I25_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_100P_1_I25_1_TQ[0]));
and2 N107P_1_100P_1_I25_1_I8_1_I6_1 (.o(N107P_1_100P_1_I25_1_I8_1_M1[0]), .i0(N107P_1_100P_1_D0), .i1(XGND));
fdce N107P_1_100P_1_I25_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[16]), .d(N107P_1_100P_1_I25_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_100P_1_I25_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_100P_1_I25_1_I13_1 (.o(N107P_1_100P_1_I25_1_L_CE), .i0(N107P_1_UN_1_CB4CLED_100P_CE), .i1(XGND));
xor2 N107P_1_100P_1_I25_1_I9_1 (.o(N107P_1_100P_1_I25_1_TQ[0]), .i0(XVDD), .i1(N107P_1_POINTER_ADDRESS[16]));
or2 N107P_1_100P_1_I22_1_I8_1_I5_1 (.o(N107P_1_100P_1_I22_1_MD[0]), .i0(N107P_1_100P_1_I22_1_I8_1_M1[0]), .i1(N107P_1_100P_1_I22_1_I8_1_M0[0]));
and2b1 N107P_1_100P_1_I22_1_I8_1_I7_1 (.o(N107P_1_100P_1_I22_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_100P_1_I22_1_TQ[0]));
and2 N107P_1_100P_1_I22_1_I8_1_I6_1 (.o(N107P_1_100P_1_I22_1_I8_1_M1[0]), .i0(N107P_1_100P_1_D3), .i1(XGND));
fdce N107P_1_100P_1_I22_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[19]), .d(N107P_1_100P_1_I22_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_100P_1_I22_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_100P_1_I22_1_I13_1 (.o(N107P_1_100P_1_I22_1_L_CE), .i0(N107P_1_UN_1_CB4CLED_100P_CE), .i1(XGND));
xor2 N107P_1_100P_1_I22_1_I9_1 (.o(N107P_1_100P_1_I22_1_TQ[0]), .i0(N107P_1_100P_1_T3), .i1(N107P_1_POINTER_ADDRESS[19]));
or2 N107P_1_100P_1_I18_1_I8_1_I5_1 (.o(N107P_1_100P_1_I18_1_MD[0]), .i0(N107P_1_100P_1_I18_1_I8_1_M1[0]), .i1(N107P_1_100P_1_I18_1_I8_1_M0[0]));
and2b1 N107P_1_100P_1_I18_1_I8_1_I7_1 (.o(N107P_1_100P_1_I18_1_I8_1_M0[0]), .i0(XGND), .i1(N107P_1_100P_1_I18_1_TQ[0]));
and2 N107P_1_100P_1_I18_1_I8_1_I6_1 (.o(N107P_1_100P_1_I18_1_I8_1_M1[0]), .i0(N107P_1_100P_1_D2), .i1(XGND));
fdce N107P_1_100P_1_I18_1_I12_1 (.q(N107P_1_POINTER_ADDRESS[18]), .d(N107P_1_100P_1_I18_1_MD[0]), .c(N107P_1_CLOCK), .ce(N107P_1_100P_1_I18_1_L_CE), .clr(XGND), .gr(RESET_n));
or2 N107P_1_100P_1_I18_1_I13_1 (.o(N107P_1_100P_1_I18_1_L_CE), .i0(N107P_1_UN_1_CB4CLED_100P_CE), .i1(XGND));
xor2 N107P_1_100P_1_I18_1_I9_1 (.o(N107P_1_100P_1_I18_1_TQ[0]), .i0(N107P_1_100P_1_T2), .i1(N107P_1_POINTER_ADDRESS[18]));
or2 N107P_1_100P_1_I29_1_I5_1 (.o(N107P_1_100P_1_T3), .i0(N107P_1_100P_1_I29_1_M1[0]), .i1(N107P_1_100P_1_I29_1_M0[0]));
and2b1 N107P_1_100P_1_I29_1_I7_1 (.o(N107P_1_100P_1_I29_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_100P_1_T3_DN));
and2 N107P_1_100P_1_I29_1_I6_1 (.o(N107P_1_100P_1_I29_1_M1[0]), .i0(N107P_1_100P_1_T3_UP), .i1(N_MEM_READ));
or2 N107P_1_100P_1_I24_1_I5_1 (.o(N107P_1_100P_1_T2), .i0(N107P_1_100P_1_I24_1_M1[0]), .i1(N107P_1_100P_1_I24_1_M0[0]));
and2b1 N107P_1_100P_1_I24_1_I7_1 (.o(N107P_1_100P_1_I24_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_100P_1_T2_DN));
and2 N107P_1_100P_1_I24_1_I6_1 (.o(N107P_1_100P_1_I24_1_M1[0]), .i0(N107P_1_100P_1_T2_UP), .i1(N_MEM_READ));
or2 N107P_1_100P_1_I23_1_I5_1 (.o(N107P_1_100P_1_TC), .i0(N107P_1_100P_1_I23_1_M1[0]), .i1(N107P_1_100P_1_I23_1_M0[0]));
and2b1 N107P_1_100P_1_I23_1_I7_1 (.o(N107P_1_100P_1_I23_1_M0[0]), .i0(N_MEM_READ), .i1(N107P_1_100P_1_TC_DN));
and2 N107P_1_100P_1_I23_1_I6_1 (.o(N107P_1_100P_1_I23_1_M1[0]), .i0(N107P_1_100P_1_TC_UP), .i1(N_MEM_READ));
and4b4 N107P_1_100P_1_I16_1 (.i3(N107P_1_POINTER_ADDRESS[17]), .i2(N107P_1_POINTER_ADDRESS[16]), .o(N107P_1_100P_1_TC_DN), .i1(N107P_1_POINTER_ADDRESS[19]), .i0(N107P_1_POINTER_ADDRESS[18]));
and3b3 N107P_1_100P_1_I21_1 (.i2(N107P_1_POINTER_ADDRESS[16]), .o(N107P_1_100P_1_T3_DN), .i1(N107P_1_POINTER_ADDRESS[18]), .i0(N107P_1_POINTER_ADDRESS[17]));
and2b2 N107P_1_100P_1_I20_1 (.o(N107P_1_100P_1_T2_DN), .i1(N107P_1_POINTER_ADDRESS[17]), .i0(N107P_1_POINTER_ADDRESS[16]));
and3 N107P_1_100P_1_I17_1 (.i2(N107P_1_POINTER_ADDRESS[16]), .o(N107P_1_100P_1_T3_UP), .i0(N107P_1_POINTER_ADDRESS[18]), .i1(N107P_1_POINTER_ADDRESS[17]));
and4 N107P_1_100P_1_I32_1 (.i2(N107P_1_POINTER_ADDRESS[17]), .i3(N107P_1_POINTER_ADDRESS[16]), .o(N107P_1_100P_1_TC_UP), .i0(N107P_1_POINTER_ADDRESS[19]), .i1(N107P_1_POINTER_ADDRESS[18]));
and2 N107P_1_100P_1_I31_1 (.o(N107P_1_100P_1_CEO), .i0(N107P_1_UN_1_CB4CLED_100P_CE), .i1(N107P_1_100P_1_TC));
and2 N107P_1_100P_1_I28_1 (.o(N107P_1_100P_1_T2_UP), .i0(N107P_1_POINTER_ADDRESS[17]), .i1(N107P_1_POINTER_ADDRESS[16]));
nor4 N107P_1_55P_1_28P_1 (.i2(N107P_1_55P_1_UN_1_NOR4_28P_I2), .i3(N107P_1_55P_1_UN_1_NOR4_28P_I3), .o(N107P_1_all_low), .i0(N107P_1_55P_1_UN_1_NOR4_28P_I0), .i1(N107P_1_55P_1_UN_1_NOR4_28P_I1));
or5 N107P_1_55P_1_25P_1 (.i4(N107P_1_POINTER_ADDRESS[4]), .i2(N107P_1_POINTER_ADDRESS[2]), .i3(N107P_1_POINTER_ADDRESS[3]), .o(N107P_1_55P_1_UN_1_NOR4_28P_I0), .i0(N107P_1_POINTER_ADDRESS[0]), .i1(N107P_1_POINTER_ADDRESS[1]));
or5 N107P_1_55P_1_24P_1 (.i4(N107P_1_POINTER_ADDRESS[19]), .i2(N107P_1_POINTER_ADDRESS[17]), .i3(N107P_1_POINTER_ADDRESS[18]), .o(N107P_1_55P_1_UN_1_NOR4_28P_I3), .i0(N107P_1_POINTER_ADDRESS[15]), .i1(N107P_1_POINTER_ADDRESS[16]));
or5 N107P_1_55P_1_26P_1 (.i4(N107P_1_POINTER_ADDRESS[14]), .i2(N107P_1_POINTER_ADDRESS[12]), .i3(N107P_1_POINTER_ADDRESS[13]), .o(N107P_1_55P_1_UN_1_NOR4_28P_I2), .i0(N107P_1_POINTER_ADDRESS[10]), .i1(N107P_1_POINTER_ADDRESS[11]));
or5 N107P_1_55P_1_23P_1 (.i4(N107P_1_POINTER_ADDRESS[9]), .i2(N107P_1_POINTER_ADDRESS[7]), .i3(N107P_1_POINTER_ADDRESS[8]), .o(N107P_1_55P_1_UN_1_NOR4_28P_I1), .i0(N107P_1_POINTER_ADDRESS[5]), .i1(N107P_1_POINTER_ADDRESS[6]));
and4 N107P_1_54P_1_2P_1 (.i2(N107P_1_54P_1_UN_1_AND4_2P_I2), .i3(N107P_1_54P_1_UN_1_AND4_2P_I3), .o(N107P_1_all_high), .i0(N107P_1_54P_1_UN_1_AND4_2P_I0), .i1(N107P_1_54P_1_UN_1_AND4_2P_I1));
and5 N107P_1_54P_1_25P_1 (.i4(N107P_1_POINTER_ADDRESS[4]), .i2(N107P_1_POINTER_ADDRESS[2]), .i3(N107P_1_POINTER_ADDRESS[3]), .o(N107P_1_54P_1_UN_1_AND4_2P_I0), .i0(N107P_1_POINTER_ADDRESS[0]), .i1(N107P_1_POINTER_ADDRESS[1]));
and5 N107P_1_54P_1_24P_1 (.i4(N107P_1_POINTER_ADDRESS[9]), .i2(N107P_1_POINTER_ADDRESS[7]), .i3(N107P_1_POINTER_ADDRESS[8]), .o(N107P_1_54P_1_UN_1_AND4_2P_I1), .i0(N107P_1_POINTER_ADDRESS[5]), .i1(N107P_1_POINTER_ADDRESS[6]));
and5 N107P_1_54P_1_26P_1 (.i4(N107P_1_POINTER_ADDRESS[19]), .i2(N107P_1_POINTER_ADDRESS[17]), .i3(N107P_1_POINTER_ADDRESS[18]), .o(N107P_1_54P_1_UN_1_AND4_2P_I3), .i0(N107P_1_POINTER_ADDRESS[15]), .i1(N107P_1_POINTER_ADDRESS[16]));
and5 N107P_1_54P_1_23P_1 (.i4(N107P_1_POINTER_ADDRESS[14]), .i2(N107P_1_POINTER_ADDRESS[12]), .i3(N107P_1_POINTER_ADDRESS[13]), .o(N107P_1_54P_1_UN_1_AND4_2P_I2), .i0(N107P_1_POINTER_ADDRESS[10]), .i1(N107P_1_POINTER_ADDRESS[11]));
inv N107P_1_97P_1_15P_1 (.i(N107P_1_97P_1_UN_1_INV_14P_O), .o(N107P_1_97P_1_UN_1_INV_15P_O));
inv N107P_1_97P_1_13P_1 (.i(N107P_1_97P_1_UN_1_INV_13P_I), .o(N107P_1_CLOCK));
inv N107P_1_97P_1_21P_1 (.i(N107P_1_97P_1_UN_1_INV_21P_I), .o(N107P_1_97P_1_UN_1_INV_20P_I));
inv N107P_1_97P_1_19P_1 (.i(N107P_1_97P_1_UN_1_INV_18P_O), .o(N107P_1_97P_1_UN_1_INV_13P_I));
inv N107P_1_97P_1_20P_1 (.i(N107P_1_97P_1_UN_1_INV_20P_I), .o(N107P_1_97P_1_UN_1_INV_14P_I));
inv N107P_1_97P_1_18P_1 (.i(N107P_1_97P_1_UN_1_INV_17P_O), .o(N107P_1_97P_1_UN_1_INV_18P_O));
inv N107P_1_97P_1_17P_1 (.i(N107P_1_97P_1_UN_1_INV_16P_O), .o(N107P_1_97P_1_UN_1_INV_17P_O));
inv N107P_1_97P_1_16P_1 (.i(N107P_1_97P_1_UN_1_INV_15P_O), .o(N107P_1_97P_1_UN_1_INV_16P_O));
inv N107P_1_97P_1_14P_1 (.i(N107P_1_97P_1_UN_1_INV_14P_I), .o(N107P_1_97P_1_UN_1_INV_14P_O));
inv N107P_1_97P_1_22P_1 (.i(N107P_1_DELAY_START), .o(N107P_1_97P_1_UN_1_INV_21P_I));
nand2 N107P_1_84P_1 (.o(N107P_1_DELAY_START), .i0(N_MEM_READ), .i1(N_MEM_WRITE));
buft N107P_1_47P_1_20 (.i(N107P_1_POINTER_ADDRESS[19]), .o(XDT[19]), .t(REG_CNTROL[2]));
buft N107P_1_47P_1_19 (.t(REG_CNTROL[2]), .o(XDT[18]), .i(N107P_1_POINTER_ADDRESS[18]));
buft N107P_1_47P_1_18 (.t(REG_CNTROL[2]), .o(XDT[17]), .i(N107P_1_POINTER_ADDRESS[17]));
buft N107P_1_47P_1_17 (.t(REG_CNTROL[2]), .o(XDT[16]), .i(N107P_1_POINTER_ADDRESS[16]));
buft N107P_1_47P_1_16 (.t(REG_CNTROL[2]), .o(XDT[15]), .i(N107P_1_POINTER_ADDRESS[15]));
buft N107P_1_47P_1_15 (.t(REG_CNTROL[2]), .o(XDT[14]), .i(N107P_1_POINTER_ADDRESS[14]));
buft N107P_1_47P_1_14 (.t(REG_CNTROL[2]), .o(XDT[13]), .i(N107P_1_POINTER_ADDRESS[13]));
buft N107P_1_47P_1_13 (.t(REG_CNTROL[2]), .o(XDT[12]), .i(N107P_1_POINTER_ADDRESS[12]));
buft N107P_1_47P_1_12 (.t(REG_CNTROL[2]), .o(XDT[11]), .i(N107P_1_POINTER_ADDRESS[11]));
buft N107P_1_47P_1_11 (.t(REG_CNTROL[2]), .o(XDT[10]), .i(N107P_1_POINTER_ADDRESS[10]));
buft N107P_1_47P_1_10 (.t(REG_CNTROL[2]), .o(XDT[9]), .i(N107P_1_POINTER_ADDRESS[9]));
buft N107P_1_47P_1_9 (.t(REG_CNTROL[2]), .o(XDT[8]), .i(N107P_1_POINTER_ADDRESS[8]));
buft N107P_1_47P_1_8 (.t(REG_CNTROL[2]), .o(XDT[7]), .i(N107P_1_POINTER_ADDRESS[7]));
buft N107P_1_47P_1_7 (.t(REG_CNTROL[2]), .o(XDT[6]), .i(N107P_1_POINTER_ADDRESS[6]));
buft N107P_1_47P_1_6 (.t(REG_CNTROL[2]), .o(XDT[5]), .i(N107P_1_POINTER_ADDRESS[5]));
buft N107P_1_47P_1_5 (.t(REG_CNTROL[2]), .o(XDT[4]), .i(N107P_1_POINTER_ADDRESS[4]));
buft N107P_1_47P_1_4 (.t(REG_CNTROL[2]), .o(XDT[3]), .i(N107P_1_POINTER_ADDRESS[3]));
buft N107P_1_47P_1_3 (.t(REG_CNTROL[2]), .o(XDT[2]), .i(N107P_1_POINTER_ADDRESS[2]));
buft N107P_1_47P_1_2 (.t(REG_CNTROL[2]), .o(XDT[1]), .i(N107P_1_POINTER_ADDRESS[1]));
buft N107P_1_47P_1_1 (.t(REG_CNTROL[2]), .o(XDT[0]), .i(N107P_1_POINTER_ADDRESS[0]));
inv N107P_1_110P_1 (.i(N107P_1_all_high), .o(WRITE_ENABLE));
inv N107P_1_109P_1 (.i(N107P_1_all_low), .o(READ_ENABLE));
gclk N96P_1 (.i(UN_1_AND2_121P_O), .o(WRITE_CU));
obuf N27P_1 (.i(UN_1_INV_119P_O), .o(BWRITE_ENABLE_n));
obuf N26P_1 (.i(UN_1_INV_120P_O), .o(BREAD_ENABLE_n));
obuf N129P_1 (.i(DOUT), .o(SDOUT));
obuf N128P_1 (.i(SM2), .o(M2));
aclk N123P_1 (.i(UN_1_ACLK_123P_I), .o(READ_CU));
and2 N122P_1 (.o(UN_1_ACLK_123P_I), .i0(N_MEM_READ), .i1(REG_CNTROL[4]));
and2 N121P_1 (.o(UN_1_AND2_121P_O), .i0(REG_CNTROL[3]), .i1(N_MEM_WRITE));
inv N120P_1 (.i(READ_ENABLE), .o(UN_1_INV_120P_O));
inv N119P_1 (.i(WRITE_ENABLE), .o(UN_1_INV_119P_O));
ibuf N61P_1_2 (.i(BXREG_ADD[1]), .o(XREG_ADD[1]));
ibuf N61P_1_1 (.o(XREG_ADD[0]), .i(BXREG_ADD[0]));
ibuf N81P_1 (.i(BMEM_WRITE_n), .o(N_MEM_WRITE));
ibuf N59P_1 (.i(BXREG_RD_n), .o(N_XREG_RD));
ibuf N58P_1 (.i(BXREG_WR_n), .o(N_XREG_WR));
ibuf N14P_1 (.i(BMEM_READ_n), .o(N_MEM_READ));
ibuf N127P_1 (.i(SDIN), .o(DIN));
ibuf N103P_1 (.i(BREAD_ADD_SEL_n), .o(N_READ_ADD_SEL));
ibuf N102P_1 (.i(BWRITE_ADD_SEL_n), .o(N_WRITE_ADD_SEL));
endmodule
`uselib

module fifo_ctrl_globals();

wire GR;
endmodule

