/* 
 *  Created:  < wittich 14/08/95>
 *  Time-stamp: <96/07/26 14:15:20 wittich>
 *  filename: /tape/snopcb/snolib_fec32/testpoint_ls/verilog_lib/verilog.v
 *  
 *  Comments: test point dummy model.
 *
 *  Modification History:
 *  ------------------------------
 *  14/08/95          Created.
 *  12/11/95          Made sizeable.  DFC.
 * 
 */ 

module TP_PAD_LS(A) ;
  input A;
  
endmodule /* TESTPOINT_LS */
   

