/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from xvmetrig3t.xcd on Fri Dec 13 11:34:41 1996 */
/* PART 3064PQ160-125 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module xvmetrig3t
(XVME_DIR, XREGWR_LA, XREGRD_LA, XMODSEL_n, XMEMSPACE_n, XMEMACK1_n, XLWORD_n, XDTACK_n, XDT_EN_n, XBRW_n, XBDS1_n, XBDS0_n, XBAM, XBA, SPARES, SDOUT, SDIN, M2, DUMMY_OUT, RDATA_n, RTRIG, RESET_n, PROGRAM_n, CCLK, PWRDWN_n);
   output XVME_DIR;
   output [31:0] XREGWR_LA;
   output [31:0] XREGRD_LA;
   output XMODSEL_n;
   output XMEMSPACE_n;
   input XMEMACK1_n;
   input XLWORD_n;
   output XDTACK_n;
   output XDT_EN_n;
   input XBRW_n;
   input XBDS1_n;
   input XBDS0_n;
   input [5:0] XBAM;
   input [31:0] XBA;
   input [3:0] SPARES;
   output SDOUT;
   input SDIN;
   output M2;
   output DUMMY_OUT;
   output RDATA_n;
   input RTRIG;
   input RESET_n;
   input PROGRAM_n;
   input CCLK;
   input PWRDWN_n;
wire [0:0] N199P_1_140P_1_D3;
wire [0:0] N199P_1_140P_1_D2;
wire [1:0] UN_1_IBUF_233P_O;
wire [31:0] REGWR_;
wire [31:0] REGRD_;
wire [5:0] BAM;
wire [31:0] BA;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/neubauer/xilinx/xvmetrig3t/verilog_lib/xvmetrig3t.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

nor3 N230P_1_26P_1 (.i0(BAM[1]), .o(N230P_1_UN_1_AND2_29P_I1), .i1(BAM[2]), .i2(BAM[4]));
nand2 N230P_1_28P_1 (.i0(N230P_1_UN_1_AND2_29P_O), .o(MEMSPACE_n), .i1(N230P_1_UN_1_INV_27P_O));
nand2 N230P_1_25P_1 (.i0(N230P_1_UN_1_AND2_29P_O), .o(REGSPACE_n), .i1(BAM[5]));
inv N230P_1_27P_1 (.i(BAM[5]), .o(N230P_1_UN_1_INV_27P_O));
and2 N230P_1_29P_1 (.i0(N230P_1_UN_1_AND2_24P_O), .o(N230P_1_UN_1_AND2_29P_O), .i1(N230P_1_UN_1_AND2_29P_I1));
and2 N230P_1_24P_1 (.i0(BAM[0]), .o(N230P_1_UN_1_AND2_24P_O), .i1(BAM[3]));
and4 N211P_1_43P_1_I30_1 (.i0(N211P_1_43P_1_PQ7), .o(N211P_1_43P_1_PQ47), .i1(N211P_1_43P_1_PQ6), .i2(N211P_1_43P_1_PQ5), .i3(N211P_1_43P_1_PQ4));
and4 N211P_1_43P_1_I28_1 (.i0(N211P_1_43P_1_PQ3), .o(N211P_1_43P_1_PQ03), .i1(N211P_1_43P_1_PQ2), .i2(N211P_1_43P_1_PQ1), .i3(N211P_1_43P_1_PQ0));
nand3b1 N211P_1_43P_1_I20_1 (.i0(REGSPACE_n), .o(N211P_1_UN_1_X74_521_40P_G), .i2(N211P_1_43P_1_PQ47), .i1(N211P_1_43P_1_PQ03));
xnor2 N211P_1_43P_1_I31_1 (.i0(BA[18]), .o(N211P_1_43P_1_PQ2), .i1(XGND));
xnor2 N211P_1_43P_1_I29_1 (.i0(XGND), .o(N211P_1_43P_1_PQ5), .i1(XGND));
xnor2 N211P_1_43P_1_I27_1 (.i0(BA[17]), .o(N211P_1_43P_1_PQ1), .i1(XGND));
xnor2 N211P_1_43P_1_I26_1 (.i0(BA[19]), .o(N211P_1_43P_1_PQ3), .i1(XGND));
xnor2 N211P_1_43P_1_I24_1 (.i0(XGND), .o(N211P_1_43P_1_PQ6), .i1(XGND));
xnor2 N211P_1_43P_1_I23_1 (.i0(XGND), .o(N211P_1_43P_1_PQ7), .i1(XGND));
xnor2 N211P_1_43P_1_I22_1 (.i0(BA[20]), .o(N211P_1_43P_1_PQ4), .i1(XGND));
xnor2 N211P_1_43P_1_I19_1 (.i0(BA[16]), .o(N211P_1_43P_1_PQ0), .i1(XGND));
and4 N211P_1_42P_1_I30_1 (.i0(N211P_1_42P_1_PQ7), .o(N211P_1_42P_1_PQ47), .i1(N211P_1_42P_1_PQ6), .i2(N211P_1_42P_1_PQ5), .i3(N211P_1_42P_1_PQ4));
and4 N211P_1_42P_1_I28_1 (.i0(N211P_1_42P_1_PQ3), .o(N211P_1_42P_1_PQ03), .i1(N211P_1_42P_1_PQ2), .i2(N211P_1_42P_1_PQ1), .i3(N211P_1_42P_1_PQ0));
nand3b1 N211P_1_42P_1_I20_1 (.i0(N211P_1_UN_1_X74_521_41P_PEQ), .o(MEMADEN_n), .i2(N211P_1_42P_1_PQ47), .i1(N211P_1_42P_1_PQ03));
xnor2 N211P_1_42P_1_I31_1 (.i0(BA[31]), .o(N211P_1_42P_1_PQ2), .i1(XGND));
xnor2 N211P_1_42P_1_I29_1 (.i0(XGND), .o(N211P_1_42P_1_PQ5), .i1(XGND));
xnor2 N211P_1_42P_1_I27_1 (.i0(BA[30]), .o(N211P_1_42P_1_PQ1), .i1(XGND));
xnor2 N211P_1_42P_1_I26_1 (.i0(XGND), .o(N211P_1_42P_1_PQ3), .i1(XGND));
xnor2 N211P_1_42P_1_I24_1 (.i0(XGND), .o(N211P_1_42P_1_PQ6), .i1(XGND));
xnor2 N211P_1_42P_1_I23_1 (.i0(XGND), .o(N211P_1_42P_1_PQ7), .i1(XGND));
xnor2 N211P_1_42P_1_I22_1 (.i0(XGND), .o(N211P_1_42P_1_PQ4), .i1(XGND));
xnor2 N211P_1_42P_1_I19_1 (.i0(BA[29]), .o(N211P_1_42P_1_PQ0), .i1(XGND));
and4 N211P_1_41P_1_I30_1 (.i0(N211P_1_41P_1_PQ7), .o(N211P_1_41P_1_PQ47), .i1(N211P_1_41P_1_PQ6), .i2(N211P_1_41P_1_PQ5), .i3(N211P_1_41P_1_PQ4));
and4 N211P_1_41P_1_I28_1 (.i0(N211P_1_41P_1_PQ3), .o(N211P_1_41P_1_PQ03), .i1(N211P_1_41P_1_PQ2), .i2(N211P_1_41P_1_PQ1), .i3(N211P_1_41P_1_PQ0));
nand3b1 N211P_1_41P_1_I20_1 (.i0(MEMSPACE_n), .o(N211P_1_UN_1_X74_521_41P_PEQ), .i2(N211P_1_41P_1_PQ47), .i1(N211P_1_41P_1_PQ03));
xnor2 N211P_1_41P_1_I31_1 (.i0(BA[23]), .o(N211P_1_41P_1_PQ2), .i1(XGND));
xnor2 N211P_1_41P_1_I29_1 (.i0(BA[26]), .o(N211P_1_41P_1_PQ5), .i1(XVDD));
xnor2 N211P_1_41P_1_I27_1 (.i0(BA[22]), .o(N211P_1_41P_1_PQ1), .i1(XGND));
xnor2 N211P_1_41P_1_I26_1 (.i0(BA[24]), .o(N211P_1_41P_1_PQ3), .i1(XGND));
xnor2 N211P_1_41P_1_I24_1 (.i0(BA[27]), .o(N211P_1_41P_1_PQ6), .i1(XGND));
xnor2 N211P_1_41P_1_I23_1 (.i0(BA[28]), .o(N211P_1_41P_1_PQ7), .i1(XGND));
xnor2 N211P_1_41P_1_I22_1 (.i0(BA[25]), .o(N211P_1_41P_1_PQ4), .i1(XGND));
xnor2 N211P_1_41P_1_I19_1 (.i0(BA[21]), .o(N211P_1_41P_1_PQ0), .i1(XGND));
and4 N211P_1_40P_1_I30_1 (.i0(N211P_1_40P_1_PQ7), .o(N211P_1_40P_1_PQ47), .i1(N211P_1_40P_1_PQ6), .i2(N211P_1_40P_1_PQ5), .i3(N211P_1_40P_1_PQ4));
and4 N211P_1_40P_1_I28_1 (.i0(N211P_1_40P_1_PQ3), .o(N211P_1_40P_1_PQ03), .i1(N211P_1_40P_1_PQ2), .i2(N211P_1_40P_1_PQ1), .i3(N211P_1_40P_1_PQ0));
nand3b1 N211P_1_40P_1_I20_1 (.i0(N211P_1_UN_1_X74_521_40P_G), .o(REGADEN_n), .i2(N211P_1_40P_1_PQ47), .i1(N211P_1_40P_1_PQ03));
xnor2 N211P_1_40P_1_I31_1 (.i0(BA[13]), .o(N211P_1_40P_1_PQ2), .i1(XVDD));
xnor2 N211P_1_40P_1_I29_1 (.i0(XGND), .o(N211P_1_40P_1_PQ5), .i1(XGND));
xnor2 N211P_1_40P_1_I27_1 (.i0(BA[12]), .o(N211P_1_40P_1_PQ1), .i1(XGND));
xnor2 N211P_1_40P_1_I26_1 (.i0(BA[14]), .o(N211P_1_40P_1_PQ3), .i1(XGND));
xnor2 N211P_1_40P_1_I24_1 (.i0(XGND), .o(N211P_1_40P_1_PQ6), .i1(XGND));
xnor2 N211P_1_40P_1_I23_1 (.i0(XGND), .o(N211P_1_40P_1_PQ7), .i1(XGND));
xnor2 N211P_1_40P_1_I22_1 (.i0(BA[15]), .o(N211P_1_40P_1_PQ4), .i1(XVDD));
xnor2 N211P_1_40P_1_I19_1 (.i0(BA[11]), .o(N211P_1_40P_1_PQ0), .i1(XGND));
nand5b4 N199P_1_190P_1_167P_1_I40_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i3(BA[5]), .o(REGWR_[16]), .i2(BA[4]), .i1(BA[3]), .i0(BA[2]));
nand5 N199P_1_190P_1_167P_1_I34_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGWR_[31]), .i1(BA[4]), .i2(BA[3]), .i3(BA[2]));
nand5b2 N199P_1_190P_1_167P_1_I39_1 (.i4(BA[3]), .i1(BA[2]), .o(REGWR_[26]), .i0(BA[4]), .i3(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_167P_1_I37_1 (.i4(BA[3]), .i1(BA[5]), .o(REGWR_[22]), .i0(BA[2]), .i3(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_167P_1_I36_1 (.i4(BA[2]), .i1(BA[5]), .o(REGWR_[21]), .i0(BA[3]), .i3(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_167P_1_I32_1 (.i4(BA[2]), .i1(BA[3]), .o(REGWR_[25]), .i0(BA[4]), .i3(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_167P_1_I31_1 (.i4(BA[4]), .i1(BA[2]), .o(REGWR_[28]), .i0(BA[3]), .i3(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_167P_1_I30_1 (.i4(BA[3]), .i1(BA[4]), .o(REGWR_[19]), .i0(BA[5]), .i3(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[2]));
nand5b3 N199P_1_190P_1_167P_1_I38_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGWR_[20]), .i1(BA[3]), .i0(BA[5]), .i3(BA[4]));
nand5b3 N199P_1_190P_1_167P_1_I35_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGWR_[24]), .i1(BA[3]), .i0(BA[4]), .i3(BA[5]));
nand5b3 N199P_1_190P_1_167P_1_I27_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[3]), .o(REGWR_[17]), .i1(BA[4]), .i0(BA[5]), .i3(BA[2]));
nand5b3 N199P_1_190P_1_167P_1_I26_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGWR_[18]), .i1(BA[5]), .i0(BA[4]), .i3(BA[3]));
nand5b1 N199P_1_190P_1_167P_1_I41_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGWR_[23]), .i3(BA[4]), .i2(BA[3]), .i1(BA[2]));
nand5b1 N199P_1_190P_1_167P_1_I33_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i0(BA[4]), .o(REGWR_[27]), .i3(BA[2]), .i2(BA[3]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_167P_1_I25_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i0(BA[2]), .o(REGWR_[30]), .i3(BA[3]), .i2(BA[4]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_167P_1_I29_1 (.i4(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i0(BA[3]), .o(REGWR_[29]), .i3(BA[2]), .i2(BA[4]), .i1(BA[5]));
nor2 N199P_1_190P_1_167P_1_I28_1 (.i0(N199P_1_WREN_n), .o(N199P_1_190P_1_167P_1_UN_1_NAND5_I34_I4), .i1(N199P_1_REG16_31_n));
nand5b4 N199P_1_190P_1_146P_1_I40_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i3(BA[5]), .o(REGWR_[0]), .i2(BA[4]), .i1(BA[3]), .i0(BA[2]));
nand5 N199P_1_190P_1_146P_1_I34_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGWR_[15]), .i1(BA[4]), .i2(BA[3]), .i3(BA[2]));
nand5b2 N199P_1_190P_1_146P_1_I39_1 (.i4(BA[3]), .i1(BA[2]), .o(REGWR_[10]), .i0(BA[4]), .i3(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_146P_1_I37_1 (.i4(BA[3]), .i1(BA[5]), .o(REGWR_[6]), .i0(BA[2]), .i3(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_146P_1_I36_1 (.i4(BA[2]), .i1(BA[5]), .o(REGWR_[5]), .i0(BA[3]), .i3(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_146P_1_I32_1 (.i4(BA[2]), .i1(BA[3]), .o(REGWR_[9]), .i0(BA[4]), .i3(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_146P_1_I31_1 (.i4(BA[4]), .i1(BA[2]), .o(REGWR_[12]), .i0(BA[3]), .i3(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_146P_1_I30_1 (.i4(BA[3]), .i1(BA[4]), .o(REGWR_[3]), .i0(BA[5]), .i3(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[2]));
nand5b3 N199P_1_190P_1_146P_1_I38_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGWR_[4]), .i1(BA[3]), .i0(BA[5]), .i3(BA[4]));
nand5b3 N199P_1_190P_1_146P_1_I35_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGWR_[8]), .i1(BA[3]), .i0(BA[4]), .i3(BA[5]));
nand5b3 N199P_1_190P_1_146P_1_I27_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[3]), .o(REGWR_[1]), .i1(BA[4]), .i0(BA[5]), .i3(BA[2]));
nand5b3 N199P_1_190P_1_146P_1_I26_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGWR_[2]), .i1(BA[5]), .i0(BA[4]), .i3(BA[3]));
nand5b1 N199P_1_190P_1_146P_1_I41_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGWR_[7]), .i3(BA[4]), .i2(BA[3]), .i1(BA[2]));
nand5b1 N199P_1_190P_1_146P_1_I33_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i0(BA[4]), .o(REGWR_[11]), .i3(BA[2]), .i2(BA[3]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_146P_1_I25_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i0(BA[2]), .o(REGWR_[14]), .i3(BA[3]), .i2(BA[4]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_146P_1_I29_1 (.i4(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i0(BA[3]), .o(REGWR_[13]), .i3(BA[2]), .i2(BA[4]), .i1(BA[5]));
nor2 N199P_1_190P_1_146P_1_I28_1 (.i0(N199P_1_WREN_n), .o(N199P_1_190P_1_146P_1_UN_1_NAND5_I34_I4), .i1(N199P_1_REG0_15_n));
nand5b4 N199P_1_190P_1_139P_1_I40_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i3(BA[5]), .o(REGRD_[0]), .i2(BA[4]), .i1(BA[3]), .i0(BA[2]));
nand5 N199P_1_190P_1_139P_1_I34_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGRD_[15]), .i1(BA[4]), .i2(BA[3]), .i3(BA[2]));
nand5b2 N199P_1_190P_1_139P_1_I39_1 (.i4(BA[3]), .i1(BA[2]), .o(REGRD_[10]), .i0(BA[4]), .i3(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_139P_1_I37_1 (.i4(BA[3]), .i1(BA[5]), .o(REGRD_[6]), .i0(BA[2]), .i3(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_139P_1_I36_1 (.i4(BA[2]), .i1(BA[5]), .o(REGRD_[5]), .i0(BA[3]), .i3(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_139P_1_I32_1 (.i4(BA[2]), .i1(BA[3]), .o(REGRD_[9]), .i0(BA[4]), .i3(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_139P_1_I31_1 (.i4(BA[4]), .i1(BA[2]), .o(REGRD_[12]), .i0(BA[3]), .i3(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_139P_1_I30_1 (.i4(BA[3]), .i1(BA[4]), .o(REGRD_[3]), .i0(BA[5]), .i3(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[2]));
nand5b3 N199P_1_190P_1_139P_1_I38_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGRD_[4]), .i1(BA[3]), .i0(BA[5]), .i3(BA[4]));
nand5b3 N199P_1_190P_1_139P_1_I35_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGRD_[8]), .i1(BA[3]), .i0(BA[4]), .i3(BA[5]));
nand5b3 N199P_1_190P_1_139P_1_I27_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[3]), .o(REGRD_[1]), .i1(BA[4]), .i0(BA[5]), .i3(BA[2]));
nand5b3 N199P_1_190P_1_139P_1_I26_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGRD_[2]), .i1(BA[5]), .i0(BA[4]), .i3(BA[3]));
nand5b1 N199P_1_190P_1_139P_1_I41_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGRD_[7]), .i3(BA[4]), .i2(BA[3]), .i1(BA[2]));
nand5b1 N199P_1_190P_1_139P_1_I33_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i0(BA[4]), .o(REGRD_[11]), .i3(BA[2]), .i2(BA[3]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_139P_1_I25_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i0(BA[2]), .o(REGRD_[14]), .i3(BA[3]), .i2(BA[4]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_139P_1_I29_1 (.i4(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i0(BA[3]), .o(REGRD_[13]), .i3(BA[2]), .i2(BA[4]), .i1(BA[5]));
nor2 N199P_1_190P_1_139P_1_I28_1 (.i0(VME_DIR), .o(N199P_1_190P_1_139P_1_UN_1_NAND5_I34_I4), .i1(N199P_1_REG0_15_n));
nand5b4 N199P_1_190P_1_138P_1_I40_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i3(BA[5]), .o(REGRD_[16]), .i2(BA[4]), .i1(BA[3]), .i0(BA[2]));
nand5 N199P_1_190P_1_138P_1_I34_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGRD_[31]), .i1(BA[4]), .i2(BA[3]), .i3(BA[2]));
nand5b2 N199P_1_190P_1_138P_1_I39_1 (.i4(BA[3]), .i1(BA[2]), .o(REGRD_[26]), .i0(BA[4]), .i3(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_138P_1_I37_1 (.i4(BA[3]), .i1(BA[5]), .o(REGRD_[22]), .i0(BA[2]), .i3(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_138P_1_I36_1 (.i4(BA[2]), .i1(BA[5]), .o(REGRD_[21]), .i0(BA[3]), .i3(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[4]));
nand5b2 N199P_1_190P_1_138P_1_I32_1 (.i4(BA[2]), .i1(BA[3]), .o(REGRD_[25]), .i0(BA[4]), .i3(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_138P_1_I31_1 (.i4(BA[4]), .i1(BA[2]), .o(REGRD_[28]), .i0(BA[3]), .i3(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[5]));
nand5b2 N199P_1_190P_1_138P_1_I30_1 (.i4(BA[3]), .i1(BA[4]), .o(REGRD_[19]), .i0(BA[5]), .i3(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[2]));
nand5b3 N199P_1_190P_1_138P_1_I38_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGRD_[20]), .i1(BA[3]), .i0(BA[5]), .i3(BA[4]));
nand5b3 N199P_1_190P_1_138P_1_I35_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGRD_[24]), .i1(BA[3]), .i0(BA[4]), .i3(BA[5]));
nand5b3 N199P_1_190P_1_138P_1_I27_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[3]), .o(REGRD_[17]), .i1(BA[4]), .i0(BA[5]), .i3(BA[2]));
nand5b3 N199P_1_190P_1_138P_1_I26_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i2(BA[2]), .o(REGRD_[18]), .i1(BA[5]), .i0(BA[4]), .i3(BA[3]));
nand5b1 N199P_1_190P_1_138P_1_I41_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i0(BA[5]), .o(REGRD_[23]), .i3(BA[4]), .i2(BA[3]), .i1(BA[2]));
nand5b1 N199P_1_190P_1_138P_1_I33_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i0(BA[4]), .o(REGRD_[27]), .i3(BA[2]), .i2(BA[3]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_138P_1_I25_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i0(BA[2]), .o(REGRD_[30]), .i3(BA[3]), .i2(BA[4]), .i1(BA[5]));
nand5b1 N199P_1_190P_1_138P_1_I29_1 (.i4(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i0(BA[3]), .o(REGRD_[29]), .i3(BA[2]), .i2(BA[4]), .i1(BA[5]));
nor2 N199P_1_190P_1_138P_1_I28_1 (.i0(VME_DIR), .o(N199P_1_190P_1_138P_1_UN_1_NAND5_I34_I4), .i1(N199P_1_REG16_31_n));
and3b1 N199P_1_140P_1_I13_1 (.i0(BA[8]), .o(N199P_1_REG16_31), .i2(BA[7]), .i1(N199P_1_UN_1_D2_4E_140P_E));
and3b1 N199P_1_140P_1_I12_1 (.i0(BA[7]), .o(N199P_1_140P_1_D2[0]), .i2(BA[8]), .i1(N199P_1_UN_1_D2_4E_140P_E));
and3b2 N199P_1_140P_1_I9_1 (.i1(BA[7]), .o(N199P_1_REG0_15), .i0(BA[8]), .i2(N199P_1_UN_1_D2_4E_140P_E));
and3 N199P_1_140P_1_I11_1 (.i0(BA[8]), .o(N199P_1_140P_1_D3[0]), .i1(BA[7]), .i2(N199P_1_UN_1_D2_4E_140P_E));
or2 N199P_1_172P_1 (.i0(REGSPACE_n), .o(N199P_1_REGSEL_n), .i1(MODSEL_n));
or2 N199P_1_171P_1 (.i0(BRW_n), .o(N199P_1_UN_1_INV_173P_I), .i1(N199P_1_REGSEL_n));
inv N199P_1_189P_1 (.i(N199P_1_REG0_15), .o(N199P_1_REG0_15_n));
inv N199P_1_188P_1 (.i(N199P_1_REG16_31), .o(N199P_1_REG16_31_n));
inv N199P_1_184P_1 (.i(BRW_n), .o(VME_DIR));
inv N199P_1_181P_1 (.i(N199P_1_UN_1_INV_181P_I), .o(N199P_1_UN_1_INV_181P_O));
inv N199P_1_169P_1 (.i(N199P_1_UN_1_INV_169P_I), .o(N199P_1_UN_1_INV_169P_O));
inv N199P_1_164P_1 (.i(N199P_1_UN_1_INV_163P_O), .o(N199P_1_UN_1_INV_164P_O));
inv N199P_1_163P_1 (.i(N199P_1_UN_1_INV_162P_O), .o(N199P_1_UN_1_INV_163P_O));
inv N199P_1_162P_1 (.i(N199P_1_UN_1_INV_161P_O), .o(N199P_1_UN_1_INV_162P_O));
inv N199P_1_161P_1 (.i(N199P_1_UN_1_INV_160P_O), .o(N199P_1_UN_1_INV_161P_O));
inv N199P_1_160P_1 (.i(N199P_1_UN_1_INV_159P_O), .o(N199P_1_UN_1_INV_160P_O));
inv N199P_1_159P_1 (.i(N199P_1_UN_1_INV_159P_I), .o(N199P_1_UN_1_INV_159P_O));
inv N199P_1_186P_1 (.i(N199P_1_UN_1_INV_181P_O), .o(N199P_1_UN_1_INV_186P_O));
inv N199P_1_182P_1 (.i(N199P_1_UN_1_INV_169P_O), .o(N199P_1_UN_1_INV_181P_I));
inv N199P_1_179P_1 (.i(N199P_1_UN_1_INV_179P_I), .o(N199P_1_UN_1_INV_178P_I));
inv N199P_1_178P_1 (.i(N199P_1_UN_1_INV_178P_I), .o(N199P_1_UN_1_INV_177P_I));
inv N199P_1_177P_1 (.i(N199P_1_UN_1_INV_177P_I), .o(N199P_1_UN_1_INV_176P_I));
inv N199P_1_176P_1 (.i(N199P_1_UN_1_INV_176P_I), .o(N199P_1_UN_1_INV_159P_I));
inv N199P_1_173P_1 (.i(N199P_1_UN_1_INV_173P_I), .o(N199P_1_UN_1_INV_169P_I));
inv N199P_1_166P_1 (.i(N199P_1_UN_1_INV_165P_O), .o(UN_1_AND2_216P_I1));
inv N199P_1_165P_1 (.i(N199P_1_UN_1_INV_164P_O), .o(N199P_1_UN_1_INV_165P_O));
nor2 N199P_1_118P_1 (.i0(N199P_1_REGSEL_n), .o(N199P_1_UN_1_D2_4E_140P_E), .i1(BA[9]));
or3 N199P_1_185P_1 (.i0(BRW_n), .o(N199P_1_WREN_n), .i1(N199P_1_UN_1_INV_186P_O), .i2(N199P_1_REGSEL_n));
and2 N199P_1_187P_1 (.i0(N199P_1_REG0_15_n), .o(N199P_1_UN_1_INV_179P_I), .i1(N199P_1_REG16_31_n));
and3 N228P_1 (.i0(BA[1]), .o(UN_1_AND3_228P_O), .i1(BA[6]), .i2(BA[10]));
or3 N225P_1 (.i0(BDS0_n), .o(UN_1_OR3_225P_O), .i1(BDS1_n), .i2(LWORD_n));
or4 N219P_1 (.i0(UN_1_OR3_225P_O), .o(MODSEL_n), .i1(UN_1_AND2_165P_O), .i2(BA[0]), .i3(UN_1_AND2_166P_O));
ibuf N198P_1_6 (.i(XBAM[5]), .o(BAM[5]));
ibuf N198P_1_5 (.o(BAM[4]), .i(XBAM[4]));
ibuf N198P_1_4 (.o(BAM[3]), .i(XBAM[3]));
ibuf N198P_1_3 (.o(BAM[2]), .i(XBAM[2]));
ibuf N198P_1_2 (.o(BAM[1]), .i(XBAM[1]));
ibuf N198P_1_1 (.o(BAM[0]), .i(XBAM[0]));
ibuf N233P_1_2 (.i(SPARES[3]), .o(UN_1_IBUF_233P_O[1]));
ibuf N233P_1_1 (.o(UN_1_IBUF_233P_O[0]), .i(SPARES[2]));
ibuf N242P_1 (.i(SDIN), .o(UN_1_IBUF_242P_O));
ibuf N224P_1 (.i(XLWORD_n), .o(LWORD_n));
ibuf N215P_1 (.i(XMEMACK1_n), .o(MEMACK1_n));
ibuf N197P_1 (.i(XBDS1_n), .o(BDS1_n));
ibuf N196P_1 (.i(XBDS0_n), .o(BDS0_n));
ibuf N195P_1 (.i(XBRW_n), .o(BRW_n));
ibuf N210P_1_32 (.i(XBA[31]), .o(BA[31]));
ibuf N210P_1_31 (.o(BA[30]), .i(XBA[30]));
ibuf N210P_1_30 (.o(BA[29]), .i(XBA[29]));
ibuf N210P_1_29 (.o(BA[28]), .i(XBA[28]));
ibuf N210P_1_28 (.o(BA[27]), .i(XBA[27]));
ibuf N210P_1_27 (.o(BA[26]), .i(XBA[26]));
ibuf N210P_1_26 (.o(BA[25]), .i(XBA[25]));
ibuf N210P_1_25 (.o(BA[24]), .i(XBA[24]));
ibuf N210P_1_24 (.o(BA[23]), .i(XBA[23]));
ibuf N210P_1_23 (.o(BA[22]), .i(XBA[22]));
ibuf N210P_1_22 (.o(BA[21]), .i(XBA[21]));
ibuf N210P_1_21 (.o(BA[20]), .i(XBA[20]));
ibuf N210P_1_20 (.o(BA[19]), .i(XBA[19]));
ibuf N210P_1_19 (.o(BA[18]), .i(XBA[18]));
ibuf N210P_1_18 (.o(BA[17]), .i(XBA[17]));
ibuf N210P_1_17 (.o(BA[16]), .i(XBA[16]));
ibuf N210P_1_16 (.o(BA[15]), .i(XBA[15]));
ibuf N210P_1_15 (.o(BA[14]), .i(XBA[14]));
ibuf N210P_1_14 (.o(BA[13]), .i(XBA[13]));
ibuf N210P_1_13 (.o(BA[12]), .i(XBA[12]));
ibuf N210P_1_12 (.o(BA[11]), .i(XBA[11]));
ibuf N210P_1_11 (.o(BA[10]), .i(XBA[10]));
ibuf N210P_1_10 (.o(BA[9]), .i(XBA[9]));
ibuf N210P_1_9 (.o(BA[8]), .i(XBA[8]));
ibuf N210P_1_8 (.o(BA[7]), .i(XBA[7]));
ibuf N210P_1_7 (.o(BA[6]), .i(XBA[6]));
ibuf N210P_1_6 (.o(BA[5]), .i(XBA[5]));
ibuf N210P_1_5 (.o(BA[4]), .i(XBA[4]));
ibuf N210P_1_4 (.o(BA[3]), .i(XBA[3]));
ibuf N210P_1_3 (.o(BA[2]), .i(XBA[2]));
ibuf N210P_1_2 (.o(BA[1]), .i(XBA[1]));
ibuf N210P_1_1 (.o(BA[0]), .i(XBA[0]));
obuf N244P_1_2 (.i(UN_1_IBUF_233P_O[1]), .o(SPARES[1]));
obuf N244P_1_1 (.o(SPARES[0]), .i(UN_1_IBUF_233P_O[0]));
obuf N241P_1 (.i(UN_1_IBUF_242P_O), .o(SDOUT));
obuf N240P_1 (.i(XVDD), .o(M2));
obuf N226P_1 (.i(UN_1_AND3_228P_O), .o(DUMMY_OUT));
obuf N217P_1 (.i(DTACK_n), .o(XDTACK_n));
obuf N180P_1 (.i(DT_EN_n), .o(XDT_EN_n));
obuf N176P_1 (.i(VME_DIR), .o(XVME_DIR));
obuf N172P_1 (.i(MODSEL_n), .o(XMODSEL_n));
obuf N171P_1 (.i(MEMSPACE_n), .o(XMEMSPACE_n));
obuf N179P_1_32 (.i(REGRD_[31]), .o(XREGRD_LA[31]));
obuf N179P_1_31 (.o(XREGRD_LA[30]), .i(REGRD_[30]));
obuf N179P_1_30 (.o(XREGRD_LA[29]), .i(REGRD_[29]));
obuf N179P_1_29 (.o(XREGRD_LA[28]), .i(REGRD_[28]));
obuf N179P_1_28 (.o(XREGRD_LA[27]), .i(REGRD_[27]));
obuf N179P_1_27 (.o(XREGRD_LA[26]), .i(REGRD_[26]));
obuf N179P_1_26 (.o(XREGRD_LA[25]), .i(REGRD_[25]));
obuf N179P_1_25 (.o(XREGRD_LA[24]), .i(REGRD_[24]));
obuf N179P_1_24 (.o(XREGRD_LA[23]), .i(REGRD_[23]));
obuf N179P_1_23 (.o(XREGRD_LA[22]), .i(REGRD_[22]));
obuf N179P_1_22 (.o(XREGRD_LA[21]), .i(REGRD_[21]));
obuf N179P_1_21 (.o(XREGRD_LA[20]), .i(REGRD_[20]));
obuf N179P_1_20 (.o(XREGRD_LA[19]), .i(REGRD_[19]));
obuf N179P_1_19 (.o(XREGRD_LA[18]), .i(REGRD_[18]));
obuf N179P_1_18 (.o(XREGRD_LA[17]), .i(REGRD_[17]));
obuf N179P_1_17 (.o(XREGRD_LA[16]), .i(REGRD_[16]));
obuf N179P_1_16 (.o(XREGRD_LA[15]), .i(REGRD_[15]));
obuf N179P_1_15 (.o(XREGRD_LA[14]), .i(REGRD_[14]));
obuf N179P_1_14 (.o(XREGRD_LA[13]), .i(REGRD_[13]));
obuf N179P_1_13 (.o(XREGRD_LA[12]), .i(REGRD_[12]));
obuf N179P_1_12 (.o(XREGRD_LA[11]), .i(REGRD_[11]));
obuf N179P_1_11 (.o(XREGRD_LA[10]), .i(REGRD_[10]));
obuf N179P_1_10 (.o(XREGRD_LA[9]), .i(REGRD_[9]));
obuf N179P_1_9 (.o(XREGRD_LA[8]), .i(REGRD_[8]));
obuf N179P_1_8 (.o(XREGRD_LA[7]), .i(REGRD_[7]));
obuf N179P_1_7 (.o(XREGRD_LA[6]), .i(REGRD_[6]));
obuf N179P_1_6 (.o(XREGRD_LA[5]), .i(REGRD_[5]));
obuf N179P_1_5 (.o(XREGRD_LA[4]), .i(REGRD_[4]));
obuf N179P_1_4 (.o(XREGRD_LA[3]), .i(REGRD_[3]));
obuf N179P_1_3 (.o(XREGRD_LA[2]), .i(REGRD_[2]));
obuf N179P_1_2 (.o(XREGRD_LA[1]), .i(REGRD_[1]));
obuf N179P_1_1 (.o(XREGRD_LA[0]), .i(REGRD_[0]));
obuf N177P_1_32 (.i(REGWR_[31]), .o(XREGWR_LA[31]));
obuf N177P_1_31 (.o(XREGWR_LA[30]), .i(REGWR_[30]));
obuf N177P_1_30 (.o(XREGWR_LA[29]), .i(REGWR_[29]));
obuf N177P_1_29 (.o(XREGWR_LA[28]), .i(REGWR_[28]));
obuf N177P_1_28 (.o(XREGWR_LA[27]), .i(REGWR_[27]));
obuf N177P_1_27 (.o(XREGWR_LA[26]), .i(REGWR_[26]));
obuf N177P_1_26 (.o(XREGWR_LA[25]), .i(REGWR_[25]));
obuf N177P_1_25 (.o(XREGWR_LA[24]), .i(REGWR_[24]));
obuf N177P_1_24 (.o(XREGWR_LA[23]), .i(REGWR_[23]));
obuf N177P_1_23 (.o(XREGWR_LA[22]), .i(REGWR_[22]));
obuf N177P_1_22 (.o(XREGWR_LA[21]), .i(REGWR_[21]));
obuf N177P_1_21 (.o(XREGWR_LA[20]), .i(REGWR_[20]));
obuf N177P_1_20 (.o(XREGWR_LA[19]), .i(REGWR_[19]));
obuf N177P_1_19 (.o(XREGWR_LA[18]), .i(REGWR_[18]));
obuf N177P_1_18 (.o(XREGWR_LA[17]), .i(REGWR_[17]));
obuf N177P_1_17 (.o(XREGWR_LA[16]), .i(REGWR_[16]));
obuf N177P_1_16 (.o(XREGWR_LA[15]), .i(REGWR_[15]));
obuf N177P_1_15 (.o(XREGWR_LA[14]), .i(REGWR_[14]));
obuf N177P_1_14 (.o(XREGWR_LA[13]), .i(REGWR_[13]));
obuf N177P_1_13 (.o(XREGWR_LA[12]), .i(REGWR_[12]));
obuf N177P_1_12 (.o(XREGWR_LA[11]), .i(REGWR_[11]));
obuf N177P_1_11 (.o(XREGWR_LA[10]), .i(REGWR_[10]));
obuf N177P_1_10 (.o(XREGWR_LA[9]), .i(REGWR_[9]));
obuf N177P_1_9 (.o(XREGWR_LA[8]), .i(REGWR_[8]));
obuf N177P_1_8 (.o(XREGWR_LA[7]), .i(REGWR_[7]));
obuf N177P_1_7 (.o(XREGWR_LA[6]), .i(REGWR_[6]));
obuf N177P_1_6 (.o(XREGWR_LA[5]), .i(REGWR_[5]));
obuf N177P_1_5 (.o(XREGWR_LA[4]), .i(REGWR_[4]));
obuf N177P_1_4 (.o(XREGWR_LA[3]), .i(REGWR_[3]));
obuf N177P_1_3 (.o(XREGWR_LA[2]), .i(REGWR_[2]));
obuf N177P_1_2 (.o(XREGWR_LA[1]), .i(REGWR_[1]));
obuf N177P_1_1 (.o(XREGWR_LA[0]), .i(REGWR_[0]));
and2 N220P_1 (.i0(DTACK_n), .o(DT_EN_n), .i1(MODSEL_n));
and2 N216P_1 (.i0(MEMACK1_n), .o(DTACK_n), .i1(UN_1_AND2_216P_I1));
and2 N166P_1 (.i0(REGADEN_n), .o(UN_1_AND2_166P_O), .i1(MEMADEN_n));
and2 N165P_1 (.i0(MEMSPACE_n), .o(UN_1_AND2_165P_O), .i1(REGSPACE_n));
endmodule
`uselib

module xvmetrig3_globals();

wire GR;
endmodule

