/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from xmemfifot.xcd on Tue Sep  3 19:36:19 1996 */
/* PART 3064PQ160-125 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module xmemfifot
(XTESTMEM2, XTESTMEM1, XSIMM_EN_, XSEL2_n, XSEL1_n, XREQ2_n, XREQ1_n, XMODSEL_n, XMEMSPACE_n, XMEMREQ2_n, XMEMACK2_n, XMEMACK1_n, XMEM_WRITE_ENABLE_n, XMDTACK, XFIFO_RESET_n, XBWR_ADD, XBRW_n, XBBA, SPARES, SDOUT, SDIN, M2, RESET_n, RDATA_n, RTRIG, PROGRAM_n, CCLK, PWRDWN_n);
   input XTESTMEM2;
   input XTESTMEM1;
   output [7:0] XSIMM_EN_;
   input XSEL2_n;
   input XSEL1_n;
   output XREQ2_n;
   output XREQ1_n;
   input XMODSEL_n;
   input XMEMSPACE_n;
   input XMEMREQ2_n;
   output XMEMACK2_n;
   output XMEMACK1_n;
   output XMEM_WRITE_ENABLE_n;
   input XMDTACK;
   input XFIFO_RESET_n;
   output [21:2] XBWR_ADD;
   input XBRW_n;
   input [24:2] XBBA;
   input [9:0] SPARES;
   output SDOUT;
   input SDIN;
   output M2;
   input RESET_n;
   output RDATA_n;
   input RTRIG;
   input PROGRAM_n;
   input CCLK;
   input PWRDWN_n;
wire [0:0] N56P_1_2P_1_I21_1_M1;
wire [0:0] N56P_1_2P_1_I21_1_M0;
wire [0:0] N56P_1_2P_1_I20_1_M1;
wire [0:0] N56P_1_2P_1_I20_1_M0;
wire [0:0] N56P_1_2P_1_I19_1_M1;
wire [0:0] N56P_1_2P_1_I19_1_M0;
wire [0:0] N56P_1_2P_1_I17_1_M1;
wire [0:0] N56P_1_2P_1_I17_1_M0;
wire [0:0] N56P_1_1P_1_I19_1_TQ;
wire [0:0] N56P_1_1P_1_I18_1_TQ;
wire [0:0] N56P_1_1P_1_I12_1_TQ;
wire [0:0] N56P_1_1P_1_I11_1_TQ;
wire [0:0] N1P_1_180P_1_77P_1_I19_1_TQ;
wire [0:0] N1P_1_180P_1_77P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_77P_1_I12_1_TQ;
wire [0:0] N1P_1_180P_1_77P_1_I11_1_TQ;
wire [0:0] N1P_1_180P_1_71P_1_I19_1_TQ;
wire [0:0] N1P_1_180P_1_71P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_71P_1_I12_1_TQ;
wire [0:0] N1P_1_180P_1_71P_1_I11_1_TQ;
wire [0:0] N1P_1_180P_1_65P_1_I19_1_TQ;
wire [0:0] N1P_1_180P_1_65P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_65P_1_I12_1_TQ;
wire [0:0] N1P_1_180P_1_65P_1_I11_1_TQ;
wire [0:0] N1P_1_180P_1_59P_1_I19_1_TQ;
wire [0:0] N1P_1_180P_1_59P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_59P_1_I12_1_TQ;
wire [0:0] N1P_1_180P_1_59P_1_I11_1_TQ;
wire [0:0] N1P_1_180P_1_53P_1_I19_1_TQ;
wire [0:0] N1P_1_180P_1_53P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_53P_1_I12_1_TQ;
wire [0:0] N1P_1_180P_1_53P_1_I11_1_TQ;
wire [0:0] N1P_1_180P_1_41P_1_I23_1_TQ;
wire [0:0] N1P_1_180P_1_41P_1_I23_1_MD;
wire [0:0] N1P_1_180P_1_41P_1_I23_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_41P_1_I23_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_41P_1_I22_1_TQ;
wire [0:0] N1P_1_180P_1_41P_1_I22_1_MD;
wire [0:0] N1P_1_180P_1_41P_1_I22_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_41P_1_I22_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_41P_1_I20_1_TQ;
wire [0:0] N1P_1_180P_1_41P_1_I20_1_MD;
wire [0:0] N1P_1_180P_1_41P_1_I20_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_41P_1_I20_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_41P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_41P_1_I18_1_MD;
wire [0:0] N1P_1_180P_1_41P_1_I18_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_41P_1_I18_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_31P_1_I23_1_TQ;
wire [0:0] N1P_1_180P_1_31P_1_I23_1_MD;
wire [0:0] N1P_1_180P_1_31P_1_I23_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_31P_1_I23_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_31P_1_I22_1_TQ;
wire [0:0] N1P_1_180P_1_31P_1_I22_1_MD;
wire [0:0] N1P_1_180P_1_31P_1_I22_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_31P_1_I22_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_31P_1_I20_1_TQ;
wire [0:0] N1P_1_180P_1_31P_1_I20_1_MD;
wire [0:0] N1P_1_180P_1_31P_1_I20_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_31P_1_I20_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_31P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_31P_1_I18_1_MD;
wire [0:0] N1P_1_180P_1_31P_1_I18_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_31P_1_I18_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_21P_1_I23_1_TQ;
wire [0:0] N1P_1_180P_1_21P_1_I23_1_MD;
wire [0:0] N1P_1_180P_1_21P_1_I23_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_21P_1_I23_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_21P_1_I22_1_TQ;
wire [0:0] N1P_1_180P_1_21P_1_I22_1_MD;
wire [0:0] N1P_1_180P_1_21P_1_I22_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_21P_1_I22_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_21P_1_I20_1_TQ;
wire [0:0] N1P_1_180P_1_21P_1_I20_1_MD;
wire [0:0] N1P_1_180P_1_21P_1_I20_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_21P_1_I20_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_21P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_21P_1_I18_1_MD;
wire [0:0] N1P_1_180P_1_21P_1_I18_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_21P_1_I18_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_11P_1_I23_1_TQ;
wire [0:0] N1P_1_180P_1_11P_1_I23_1_MD;
wire [0:0] N1P_1_180P_1_11P_1_I23_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_11P_1_I23_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_11P_1_I22_1_TQ;
wire [0:0] N1P_1_180P_1_11P_1_I22_1_MD;
wire [0:0] N1P_1_180P_1_11P_1_I22_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_11P_1_I22_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_11P_1_I20_1_TQ;
wire [0:0] N1P_1_180P_1_11P_1_I20_1_MD;
wire [0:0] N1P_1_180P_1_11P_1_I20_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_11P_1_I20_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_11P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_11P_1_I18_1_MD;
wire [0:0] N1P_1_180P_1_11P_1_I18_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_11P_1_I18_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_1P_1_I23_1_TQ;
wire [0:0] N1P_1_180P_1_1P_1_I23_1_MD;
wire [0:0] N1P_1_180P_1_1P_1_I23_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_1P_1_I23_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_1P_1_I22_1_TQ;
wire [0:0] N1P_1_180P_1_1P_1_I22_1_MD;
wire [0:0] N1P_1_180P_1_1P_1_I22_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_1P_1_I22_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_1P_1_I20_1_TQ;
wire [0:0] N1P_1_180P_1_1P_1_I20_1_MD;
wire [0:0] N1P_1_180P_1_1P_1_I20_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_1P_1_I20_1_I8_1_M0;
wire [0:0] N1P_1_180P_1_1P_1_I18_1_TQ;
wire [0:0] N1P_1_180P_1_1P_1_I18_1_MD;
wire [0:0] N1P_1_180P_1_1P_1_I18_1_I8_1_M1;
wire [0:0] N1P_1_180P_1_1P_1_I18_1_I8_1_M0;
wire [0:0] N1P_1_179P_1_74P_1_AB3;
wire [0:0] N1P_1_179P_1_74P_1_AB2;
wire [0:0] N1P_1_179P_1_74P_1_AB1;
wire [0:0] N1P_1_179P_1_74P_1_AB0;
wire [0:0] N1P_1_179P_1_70P_1_AB3;
wire [0:0] N1P_1_179P_1_70P_1_AB2;
wire [0:0] N1P_1_179P_1_70P_1_AB1;
wire [0:0] N1P_1_179P_1_70P_1_AB0;
wire [0:0] N1P_1_179P_1_66P_1_AB3;
wire [0:0] N1P_1_179P_1_66P_1_AB2;
wire [0:0] N1P_1_179P_1_66P_1_AB1;
wire [0:0] N1P_1_179P_1_66P_1_AB0;
wire [0:0] N1P_1_179P_1_62P_1_AB3;
wire [0:0] N1P_1_179P_1_62P_1_AB2;
wire [0:0] N1P_1_179P_1_62P_1_AB1;
wire [0:0] N1P_1_179P_1_62P_1_AB0;
wire [0:0] N1P_1_179P_1_58P_1_AB3;
wire [0:0] N1P_1_179P_1_58P_1_AB2;
wire [0:0] N1P_1_179P_1_58P_1_AB1;
wire [0:0] N1P_1_179P_1_58P_1_AB0;
wire [19:0] N1P_1_NEXT_READ;
wire [19:0] N1P_1_LAST_WRITE;
wire [19:0] N1P_1_LAST_READ;
wire [4:0] UN_1_IBUF_82P_O;
wire [7:0] SIMM_EN_;
wire [21:2] BWR_ADD;
wire [24:2] BBA;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/neubauer/xilinx/xmemfifot/verilog_lib/xmemfifot.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

fdce N65P_1_I8_1 (.q(UN_1_FDC_65P_Q), .d(XVDD), .c(UN_1_FDC_65P_C), .clr(UN_1_FDC_65P_CLR), .ce(XVDD), .gr(RESET_n));
nand4b3 N56P_1_6P_1_I23_1 (.i2(N56P_1_LY1), .i3(N56P_1_6P_1_E), .o(SIMM_EN_[0]), .i1(N56P_1_LY2), .i0(N56P_1_LY3));
nand4b2 N56P_1_6P_1_I25_1 (.i3(N56P_1_LY2), .i2(N56P_1_6P_1_E), .o(SIMM_EN_[2]), .i1(N56P_1_LY1), .i0(N56P_1_LY3));
nand4b2 N56P_1_6P_1_I21_1 (.i3(N56P_1_LY1), .i2(N56P_1_6P_1_E), .o(SIMM_EN_[1]), .i1(N56P_1_LY2), .i0(N56P_1_LY3));
nand4b2 N56P_1_6P_1_I20_1 (.i3(N56P_1_LY3), .i2(N56P_1_6P_1_E), .o(SIMM_EN_[4]), .i1(N56P_1_LY1), .i0(N56P_1_LY2));
nand4 N56P_1_6P_1_I17_1 (.i2(N56P_1_LY1), .i3(N56P_1_6P_1_E), .o(SIMM_EN_[7]), .i1(N56P_1_LY2), .i0(N56P_1_LY3));
and3b2 N56P_1_6P_1_I16_1 (.i2(REQ1), .o(N56P_1_6P_1_E), .i1(XGND), .i0(XGND));
nand4b1 N56P_1_6P_1_I22_1 (.i3(N56P_1_LY1), .i2(N56P_1_6P_1_E), .o(SIMM_EN_[5]), .i1(N56P_1_LY3), .i0(N56P_1_LY2));
nand4b1 N56P_1_6P_1_I15_1 (.i3(N56P_1_LY2), .i2(N56P_1_6P_1_E), .o(SIMM_EN_[6]), .i1(N56P_1_LY3), .i0(N56P_1_LY1));
nand4b1 N56P_1_6P_1_I18_1 (.i3(N56P_1_LY2), .i2(N56P_1_6P_1_E), .o(SIMM_EN_[3]), .i1(N56P_1_LY1), .i0(N56P_1_LY3));
and3b1 N56P_1_2P_1_I21_1_I6_1 (.i2(N56P_1_UN_1_CB4CE_1P_Q2), .o(N56P_1_2P_1_I21_1_M0[0]), .i1(N56P_1_2P_1_E), .i0(TESTMEM1));
and3 N56P_1_2P_1_I21_1_I10_1 (.i2(TESTMEM1), .o(N56P_1_2P_1_I21_1_M1[0]), .i1(N56P_1_2P_1_E), .i0(BBA[24]));
or2 N56P_1_2P_1_I21_1_I8_1 (.o(N56P_1_Y3), .i1(N56P_1_2P_1_I21_1_M0[0]), .i0(N56P_1_2P_1_I21_1_M1[0]));
and3b1 N56P_1_2P_1_I20_1_I6_1 (.i2(N56P_1_UN_1_CB4CE_1P_Q0), .o(N56P_1_2P_1_I20_1_M0[0]), .i1(N56P_1_2P_1_E), .i0(TESTMEM1));
and3 N56P_1_2P_1_I20_1_I10_1 (.i2(TESTMEM1), .o(N56P_1_2P_1_I20_1_M1[0]), .i1(N56P_1_2P_1_E), .i0(BBA[22]));
or2 N56P_1_2P_1_I20_1_I8_1 (.o(N56P_1_Y1), .i1(N56P_1_2P_1_I20_1_M0[0]), .i0(N56P_1_2P_1_I20_1_M1[0]));
and3b1 N56P_1_2P_1_I17_1_I6_1 (.i2(XGND), .o(N56P_1_2P_1_I17_1_M0[0]), .i1(N56P_1_2P_1_E), .i0(TESTMEM1));
and3 N56P_1_2P_1_I17_1_I10_1 (.i2(TESTMEM1), .o(N56P_1_2P_1_I17_1_M1[0]), .i1(N56P_1_2P_1_E), .i0(XGND));
or2 N56P_1_2P_1_I17_1_I8_1 (.o(N56P_1_2P_1_Y4), .i1(N56P_1_2P_1_I17_1_M0[0]), .i0(N56P_1_2P_1_I17_1_M1[0]));
and3b1 N56P_1_2P_1_I19_1_I6_1 (.i2(N56P_1_UN_1_CB4CE_1P_Q1), .o(N56P_1_2P_1_I19_1_M0[0]), .i1(N56P_1_2P_1_E), .i0(TESTMEM1));
and3 N56P_1_2P_1_I19_1_I10_1 (.i2(TESTMEM1), .o(N56P_1_2P_1_I19_1_M1[0]), .i1(N56P_1_2P_1_E), .i0(BBA[23]));
or2 N56P_1_2P_1_I19_1_I8_1 (.o(N56P_1_Y2), .i1(N56P_1_2P_1_I19_1_M0[0]), .i0(N56P_1_2P_1_I19_1_M1[0]));
inv N56P_1_2P_1_I18_1 (.i(XGND), .o(N56P_1_2P_1_E));
xor2 N56P_1_1P_1_I19_1_I8_1 (.o(N56P_1_1P_1_I19_1_TQ[0]), .i1(N56P_1_UN_1_CB4CE_1P_Q2), .i0(N56P_1_1P_1_T2));
fdce N56P_1_1P_1_I19_1_I7_1 (.q(N56P_1_UN_1_CB4CE_1P_Q2), .d(N56P_1_1P_1_I19_1_TQ[0]), .c(MEMACK1_n), .clr(N56P_1_UN_1_CB4CE_1P_CLR), .ce(XVDD), .gr(RESET_n));
xor2 N56P_1_1P_1_I18_1_I8_1 (.o(N56P_1_1P_1_I18_1_TQ[0]), .i1(N56P_1_UN_1_CB4CE_1P_Q1), .i0(N56P_1_UN_1_CB4CE_1P_Q0));
fdce N56P_1_1P_1_I18_1_I7_1 (.q(N56P_1_UN_1_CB4CE_1P_Q1), .d(N56P_1_1P_1_I18_1_TQ[0]), .c(MEMACK1_n), .clr(N56P_1_UN_1_CB4CE_1P_CLR), .ce(XVDD), .gr(RESET_n));
xor2 N56P_1_1P_1_I12_1_I8_1 (.o(N56P_1_1P_1_I12_1_TQ[0]), .i1(N56P_1_UN_1_CB4CE_1P_Q0), .i0(XVDD));
fdce N56P_1_1P_1_I12_1_I7_1 (.q(N56P_1_UN_1_CB4CE_1P_Q0), .d(N56P_1_1P_1_I12_1_TQ[0]), .c(MEMACK1_n), .clr(N56P_1_UN_1_CB4CE_1P_CLR), .ce(XVDD), .gr(RESET_n));
xor2 N56P_1_1P_1_I11_1_I8_1 (.o(N56P_1_1P_1_I11_1_TQ[0]), .i1(N56P_1_1P_1_Q3), .i0(N56P_1_1P_1_T3));
fdce N56P_1_1P_1_I11_1_I7_1 (.gr(XVDD), .q(N56P_1_1P_1_Q3), .d(N56P_1_1P_1_I11_1_TQ[0]), .c(MEMACK1_n), .clr(N56P_1_UN_1_CB4CE_1P_CLR), .ce(XVDD));
and3 N56P_1_1P_1_I13_1 (.i2(N56P_1_UN_1_CB4CE_1P_Q0), .o(N56P_1_1P_1_T3), .i1(N56P_1_UN_1_CB4CE_1P_Q1), .i0(N56P_1_UN_1_CB4CE_1P_Q2));
and4 N56P_1_1P_1_I10_1 (.i2(N56P_1_UN_1_CB4CE_1P_Q1), .i3(N56P_1_UN_1_CB4CE_1P_Q0), .o(N56P_1_1P_1_TC), .i1(N56P_1_UN_1_CB4CE_1P_Q2), .i0(N56P_1_1P_1_Q3));
and2 N56P_1_1P_1_I16_1 (.o(N56P_1_1P_1_CEO), .i1(N56P_1_1P_1_TC), .i0(XVDD));
and2 N56P_1_1P_1_I14_1 (.o(N56P_1_1P_1_T2), .i1(N56P_1_UN_1_CB4CE_1P_Q0), .i0(N56P_1_UN_1_CB4CE_1P_Q1));
fdce N56P_1_3P_1_I6_1 (.q(N56P_1_LY2), .d(N56P_1_Y2), .c(MEMREQ1), .clr(XGND), .ce(XVDD), .gr(RESET_n));
fdce N56P_1_5P_1_I6_1 (.q(N56P_1_LY1), .d(N56P_1_Y1), .c(MEMREQ1), .clr(XGND), .ce(XVDD), .gr(RESET_n));
fdce N56P_1_7P_1_I6_1 (.q(N56P_1_LY3), .d(N56P_1_Y3), .c(MEMREQ1), .clr(XGND), .ce(XVDD), .gr(RESET_n));
inv N56P_1_27P_1 (.i(READ_BLKACK_n), .o(N56P_1_UN_1_CB4CE_1P_CLR));
fdce N42P_1_25P_1_I8_1 (.q(N42P_1_REQ2_OUT), .d(XVDD), .c(N42P_1_REQ2_CLK), .clr(N42P_1_REQ2_CLR), .ce(XVDD), .gr(RESET_n));
fdce N42P_1_24P_1_I8_1 (.q(N42P_1_UN_1_FDC_24P_Q), .d(XVDD), .c(N42P_1_MDTACK_n), .clr(N42P_1_STILL_REQ_n), .ce(XVDD), .gr(RESET_n));
nand2 N42P_1_13P_1 (.o(N42P_1_STILL_REQ_n), .i1(N42P_1_REQ2_IN), .i0(REQ2_n));
and2 N42P_1_23P_1 (.o(N42P_1_REQ2_CLK), .i1(N42P_1_REQ2_IN), .i0(N42P_1_STILL_REQ_CLK));
nor2 N42P_1_22P_1 (.o(N42P_1_REQ2_CLR), .i1(N42P_1_MDTACK_n), .i0(REQ2_n));
or2 N42P_1_19P_1 (.o(N42P_1_STILL_REQ_CLK), .i1(N42P_1_UN_1_FDC_24P_Q), .i0(N42P_1_MDTACK_n));
inv N42P_1_20P_1 (.i(N42P_1_REQ2_OUT), .o(REQ2_n));
inv N42P_1_18P_1 (.i(REQ2_IN_n), .o(N42P_1_REQ2_IN));
inv N42P_1_17P_1 (.i(MDTACK), .o(N42P_1_MDTACK_n));
fdce N1P_1_182P_1_I8_1_20 (.q(N1P_1_LAST_WRITE[19]), .d(BWR_ADD[21]), .c(N1P_1_SEL2), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_19 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[20]), .q(N1P_1_LAST_WRITE[18]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_18 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[19]), .q(N1P_1_LAST_WRITE[17]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_17 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[18]), .q(N1P_1_LAST_WRITE[16]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_16 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[17]), .q(N1P_1_LAST_WRITE[15]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_15 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[16]), .q(N1P_1_LAST_WRITE[14]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_14 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[15]), .q(N1P_1_LAST_WRITE[13]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_13 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[14]), .q(N1P_1_LAST_WRITE[12]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_12 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[13]), .q(N1P_1_LAST_WRITE[11]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_11 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[12]), .q(N1P_1_LAST_WRITE[10]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_10 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[11]), .q(N1P_1_LAST_WRITE[9]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_9 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[10]), .q(N1P_1_LAST_WRITE[8]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_8 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[9]), .q(N1P_1_LAST_WRITE[7]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_7 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[8]), .q(N1P_1_LAST_WRITE[6]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_6 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[7]), .q(N1P_1_LAST_WRITE[5]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_5 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[6]), .q(N1P_1_LAST_WRITE[4]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_4 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[5]), .q(N1P_1_LAST_WRITE[3]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_3 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[4]), .q(N1P_1_LAST_WRITE[2]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_2 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[3]), .q(N1P_1_LAST_WRITE[1]), .gr(RESET_n));
fdce N1P_1_182P_1_I8_1_1 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL2), .d(BWR_ADD[2]), .q(N1P_1_LAST_WRITE[0]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_20 (.q(N1P_1_LAST_READ[19]), .d(BBA[21]), .c(N1P_1_SEL1), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_19 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[20]), .q(N1P_1_LAST_READ[18]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_18 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[19]), .q(N1P_1_LAST_READ[17]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_17 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[18]), .q(N1P_1_LAST_READ[16]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_16 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[17]), .q(N1P_1_LAST_READ[15]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_15 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[16]), .q(N1P_1_LAST_READ[14]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_14 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[15]), .q(N1P_1_LAST_READ[13]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_13 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[14]), .q(N1P_1_LAST_READ[12]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_12 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[13]), .q(N1P_1_LAST_READ[11]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_11 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[12]), .q(N1P_1_LAST_READ[10]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_10 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[11]), .q(N1P_1_LAST_READ[9]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_9 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[10]), .q(N1P_1_LAST_READ[8]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_8 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[9]), .q(N1P_1_LAST_READ[7]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_7 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[8]), .q(N1P_1_LAST_READ[6]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_6 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[7]), .q(N1P_1_LAST_READ[5]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_5 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[6]), .q(N1P_1_LAST_READ[4]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_4 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[5]), .q(N1P_1_LAST_READ[3]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_3 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[4]), .q(N1P_1_LAST_READ[2]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_2 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[3]), .q(N1P_1_LAST_READ[1]), .gr(RESET_n));
fdce N1P_1_174P_1_I8_1_1 (.ce(XVDD), .clr(N1P_1_FIFO_RESET), .c(N1P_1_SEL1), .d(BBA[2]), .q(N1P_1_LAST_READ[0]), .gr(RESET_n));
and2b1 N1P_1_180P_1_31P_1_I23_1_I8_1_I7_1 (.o(N1P_1_180P_1_31P_1_I23_1_I8_1_M0[0]), .i1(N1P_1_180P_1_31P_1_I23_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_31P_1_I23_1_I8_1_I6_1 (.o(N1P_1_180P_1_31P_1_I23_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[7]));
or2 N1P_1_180P_1_31P_1_I23_1_I8_1_I5_1 (.o(N1P_1_180P_1_31P_1_I23_1_MD[0]), .i1(N1P_1_180P_1_31P_1_I23_1_I8_1_M0[0]), .i0(N1P_1_180P_1_31P_1_I23_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_31P_1_I23_1_I9_1 (.o(N1P_1_180P_1_31P_1_I23_1_TQ[0]), .i1(N1P_1_NEXT_READ[5]), .i0(N1P_1_NEXT_READ[4]));
fdce N1P_1_180P_1_31P_1_I23_1_I12_1 (.q(N1P_1_NEXT_READ[5]), .d(N1P_1_180P_1_31P_1_I23_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_31P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_31P_1_I23_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_31P_1_I23_1_I13_1 (.o(N1P_1_180P_1_31P_1_I23_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_31P_1_I22_1_I8_1_I7_1 (.o(N1P_1_180P_1_31P_1_I22_1_I8_1_M0[0]), .i1(N1P_1_180P_1_31P_1_I22_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_31P_1_I22_1_I8_1_I6_1 (.o(N1P_1_180P_1_31P_1_I22_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[6]));
or2 N1P_1_180P_1_31P_1_I22_1_I8_1_I5_1 (.o(N1P_1_180P_1_31P_1_I22_1_MD[0]), .i1(N1P_1_180P_1_31P_1_I22_1_I8_1_M0[0]), .i0(N1P_1_180P_1_31P_1_I22_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_31P_1_I22_1_I9_1 (.o(N1P_1_180P_1_31P_1_I22_1_TQ[0]), .i1(N1P_1_NEXT_READ[4]), .i0(XVDD));
fdce N1P_1_180P_1_31P_1_I22_1_I12_1 (.q(N1P_1_NEXT_READ[4]), .d(N1P_1_180P_1_31P_1_I22_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_31P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_31P_1_I22_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_31P_1_I22_1_I13_1 (.o(N1P_1_180P_1_31P_1_I22_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_31P_1_I20_1_I8_1_I7_1 (.o(N1P_1_180P_1_31P_1_I20_1_I8_1_M0[0]), .i1(N1P_1_180P_1_31P_1_I20_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_31P_1_I20_1_I8_1_I6_1 (.o(N1P_1_180P_1_31P_1_I20_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[9]));
or2 N1P_1_180P_1_31P_1_I20_1_I8_1_I5_1 (.o(N1P_1_180P_1_31P_1_I20_1_MD[0]), .i1(N1P_1_180P_1_31P_1_I20_1_I8_1_M0[0]), .i0(N1P_1_180P_1_31P_1_I20_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_31P_1_I20_1_I9_1 (.o(N1P_1_180P_1_31P_1_I20_1_TQ[0]), .i1(N1P_1_NEXT_READ[7]), .i0(N1P_1_180P_1_31P_1_T3));
fdce N1P_1_180P_1_31P_1_I20_1_I12_1 (.q(N1P_1_NEXT_READ[7]), .d(N1P_1_180P_1_31P_1_I20_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_31P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_31P_1_I20_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_31P_1_I20_1_I13_1 (.o(N1P_1_180P_1_31P_1_I20_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_31P_1_I18_1_I8_1_I7_1 (.o(N1P_1_180P_1_31P_1_I18_1_I8_1_M0[0]), .i1(N1P_1_180P_1_31P_1_I18_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_31P_1_I18_1_I8_1_I6_1 (.o(N1P_1_180P_1_31P_1_I18_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[8]));
or2 N1P_1_180P_1_31P_1_I18_1_I8_1_I5_1 (.o(N1P_1_180P_1_31P_1_I18_1_MD[0]), .i1(N1P_1_180P_1_31P_1_I18_1_I8_1_M0[0]), .i0(N1P_1_180P_1_31P_1_I18_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_31P_1_I18_1_I9_1 (.o(N1P_1_180P_1_31P_1_I18_1_TQ[0]), .i1(N1P_1_NEXT_READ[6]), .i0(N1P_1_180P_1_31P_1_T2));
fdce N1P_1_180P_1_31P_1_I18_1_I12_1 (.q(N1P_1_NEXT_READ[6]), .d(N1P_1_180P_1_31P_1_I18_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_31P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_31P_1_I18_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_31P_1_I18_1_I13_1 (.o(N1P_1_180P_1_31P_1_I18_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and3 N1P_1_180P_1_31P_1_I21_1 (.i2(N1P_1_NEXT_READ[4]), .o(N1P_1_180P_1_31P_1_T3), .i1(N1P_1_NEXT_READ[5]), .i0(N1P_1_NEXT_READ[6]));
and4 N1P_1_180P_1_31P_1_I19_1 (.i2(N1P_1_NEXT_READ[6]), .i3(N1P_1_NEXT_READ[7]), .o(N1P_1_180P_1_UN_1_CB4CLE_31P_TC), .i1(N1P_1_NEXT_READ[5]), .i0(N1P_1_NEXT_READ[4]));
and2 N1P_1_180P_1_31P_1_I24_1 (.o(N1P_1_180P_1_31P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CLE_31P_TC), .i0(XVDD));
and2 N1P_1_180P_1_31P_1_I17_1 (.o(N1P_1_180P_1_31P_1_T2), .i1(N1P_1_NEXT_READ[4]), .i0(N1P_1_NEXT_READ[5]));
and2b1 N1P_1_180P_1_41P_1_I23_1_I8_1_I7_1 (.o(N1P_1_180P_1_41P_1_I23_1_I8_1_M0[0]), .i1(N1P_1_180P_1_41P_1_I23_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_41P_1_I23_1_I8_1_I6_1 (.o(N1P_1_180P_1_41P_1_I23_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[3]));
or2 N1P_1_180P_1_41P_1_I23_1_I8_1_I5_1 (.o(N1P_1_180P_1_41P_1_I23_1_MD[0]), .i1(N1P_1_180P_1_41P_1_I23_1_I8_1_M0[0]), .i0(N1P_1_180P_1_41P_1_I23_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_41P_1_I23_1_I9_1 (.o(N1P_1_180P_1_41P_1_I23_1_TQ[0]), .i1(N1P_1_NEXT_READ[1]), .i0(N1P_1_NEXT_READ[0]));
fdce N1P_1_180P_1_41P_1_I23_1_I12_1 (.q(N1P_1_NEXT_READ[1]), .d(N1P_1_180P_1_41P_1_I23_1_MD[0]), .c(READ_BLKACK_n), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_41P_1_I23_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_41P_1_I23_1_I13_1 (.o(N1P_1_180P_1_41P_1_I23_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_41P_1_I22_1_I8_1_I7_1 (.o(N1P_1_180P_1_41P_1_I22_1_I8_1_M0[0]), .i1(N1P_1_180P_1_41P_1_I22_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_41P_1_I22_1_I8_1_I6_1 (.o(N1P_1_180P_1_41P_1_I22_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[2]));
or2 N1P_1_180P_1_41P_1_I22_1_I8_1_I5_1 (.o(N1P_1_180P_1_41P_1_I22_1_MD[0]), .i1(N1P_1_180P_1_41P_1_I22_1_I8_1_M0[0]), .i0(N1P_1_180P_1_41P_1_I22_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_41P_1_I22_1_I9_1 (.o(N1P_1_180P_1_41P_1_I22_1_TQ[0]), .i1(N1P_1_NEXT_READ[0]), .i0(XVDD));
fdce N1P_1_180P_1_41P_1_I22_1_I12_1 (.q(N1P_1_NEXT_READ[0]), .d(N1P_1_180P_1_41P_1_I22_1_MD[0]), .c(READ_BLKACK_n), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_41P_1_I22_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_41P_1_I22_1_I13_1 (.o(N1P_1_180P_1_41P_1_I22_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_41P_1_I20_1_I8_1_I7_1 (.o(N1P_1_180P_1_41P_1_I20_1_I8_1_M0[0]), .i1(N1P_1_180P_1_41P_1_I20_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_41P_1_I20_1_I8_1_I6_1 (.o(N1P_1_180P_1_41P_1_I20_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[5]));
or2 N1P_1_180P_1_41P_1_I20_1_I8_1_I5_1 (.o(N1P_1_180P_1_41P_1_I20_1_MD[0]), .i1(N1P_1_180P_1_41P_1_I20_1_I8_1_M0[0]), .i0(N1P_1_180P_1_41P_1_I20_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_41P_1_I20_1_I9_1 (.o(N1P_1_180P_1_41P_1_I20_1_TQ[0]), .i1(N1P_1_NEXT_READ[3]), .i0(N1P_1_180P_1_41P_1_T3));
fdce N1P_1_180P_1_41P_1_I20_1_I12_1 (.q(N1P_1_NEXT_READ[3]), .d(N1P_1_180P_1_41P_1_I20_1_MD[0]), .c(READ_BLKACK_n), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_41P_1_I20_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_41P_1_I20_1_I13_1 (.o(N1P_1_180P_1_41P_1_I20_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_41P_1_I18_1_I8_1_I7_1 (.o(N1P_1_180P_1_41P_1_I18_1_I8_1_M0[0]), .i1(N1P_1_180P_1_41P_1_I18_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_41P_1_I18_1_I8_1_I6_1 (.o(N1P_1_180P_1_41P_1_I18_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[4]));
or2 N1P_1_180P_1_41P_1_I18_1_I8_1_I5_1 (.o(N1P_1_180P_1_41P_1_I18_1_MD[0]), .i1(N1P_1_180P_1_41P_1_I18_1_I8_1_M0[0]), .i0(N1P_1_180P_1_41P_1_I18_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_41P_1_I18_1_I9_1 (.o(N1P_1_180P_1_41P_1_I18_1_TQ[0]), .i1(N1P_1_NEXT_READ[2]), .i0(N1P_1_180P_1_41P_1_T2));
fdce N1P_1_180P_1_41P_1_I18_1_I12_1 (.q(N1P_1_NEXT_READ[2]), .d(N1P_1_180P_1_41P_1_I18_1_MD[0]), .c(READ_BLKACK_n), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_41P_1_I18_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_41P_1_I18_1_I13_1 (.o(N1P_1_180P_1_41P_1_I18_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and3 N1P_1_180P_1_41P_1_I21_1 (.i2(N1P_1_NEXT_READ[0]), .o(N1P_1_180P_1_41P_1_T3), .i1(N1P_1_NEXT_READ[1]), .i0(N1P_1_NEXT_READ[2]));
and4 N1P_1_180P_1_41P_1_I19_1 (.i2(N1P_1_NEXT_READ[2]), .i3(N1P_1_NEXT_READ[3]), .o(N1P_1_180P_1_UN_1_CB4CLE_41P_TC), .i1(N1P_1_NEXT_READ[1]), .i0(N1P_1_NEXT_READ[0]));
and2 N1P_1_180P_1_41P_1_I24_1 (.o(N1P_1_180P_1_41P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CLE_41P_TC), .i0(XVDD));
and2 N1P_1_180P_1_41P_1_I17_1 (.o(N1P_1_180P_1_41P_1_T2), .i1(N1P_1_NEXT_READ[0]), .i0(N1P_1_NEXT_READ[1]));
and2b1 N1P_1_180P_1_21P_1_I23_1_I8_1_I7_1 (.o(N1P_1_180P_1_21P_1_I23_1_I8_1_M0[0]), .i1(N1P_1_180P_1_21P_1_I23_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_21P_1_I23_1_I8_1_I6_1 (.o(N1P_1_180P_1_21P_1_I23_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[11]));
or2 N1P_1_180P_1_21P_1_I23_1_I8_1_I5_1 (.o(N1P_1_180P_1_21P_1_I23_1_MD[0]), .i1(N1P_1_180P_1_21P_1_I23_1_I8_1_M0[0]), .i0(N1P_1_180P_1_21P_1_I23_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_21P_1_I23_1_I9_1 (.o(N1P_1_180P_1_21P_1_I23_1_TQ[0]), .i1(N1P_1_NEXT_READ[9]), .i0(N1P_1_NEXT_READ[8]));
fdce N1P_1_180P_1_21P_1_I23_1_I12_1 (.q(N1P_1_NEXT_READ[9]), .d(N1P_1_180P_1_21P_1_I23_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_21P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_21P_1_I23_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_21P_1_I23_1_I13_1 (.o(N1P_1_180P_1_21P_1_I23_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_21P_1_I22_1_I8_1_I7_1 (.o(N1P_1_180P_1_21P_1_I22_1_I8_1_M0[0]), .i1(N1P_1_180P_1_21P_1_I22_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_21P_1_I22_1_I8_1_I6_1 (.o(N1P_1_180P_1_21P_1_I22_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[10]));
or2 N1P_1_180P_1_21P_1_I22_1_I8_1_I5_1 (.o(N1P_1_180P_1_21P_1_I22_1_MD[0]), .i1(N1P_1_180P_1_21P_1_I22_1_I8_1_M0[0]), .i0(N1P_1_180P_1_21P_1_I22_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_21P_1_I22_1_I9_1 (.o(N1P_1_180P_1_21P_1_I22_1_TQ[0]), .i1(N1P_1_NEXT_READ[8]), .i0(XVDD));
fdce N1P_1_180P_1_21P_1_I22_1_I12_1 (.q(N1P_1_NEXT_READ[8]), .d(N1P_1_180P_1_21P_1_I22_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_21P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_21P_1_I22_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_21P_1_I22_1_I13_1 (.o(N1P_1_180P_1_21P_1_I22_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_21P_1_I20_1_I8_1_I7_1 (.o(N1P_1_180P_1_21P_1_I20_1_I8_1_M0[0]), .i1(N1P_1_180P_1_21P_1_I20_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_21P_1_I20_1_I8_1_I6_1 (.o(N1P_1_180P_1_21P_1_I20_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[13]));
or2 N1P_1_180P_1_21P_1_I20_1_I8_1_I5_1 (.o(N1P_1_180P_1_21P_1_I20_1_MD[0]), .i1(N1P_1_180P_1_21P_1_I20_1_I8_1_M0[0]), .i0(N1P_1_180P_1_21P_1_I20_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_21P_1_I20_1_I9_1 (.o(N1P_1_180P_1_21P_1_I20_1_TQ[0]), .i1(N1P_1_NEXT_READ[11]), .i0(N1P_1_180P_1_21P_1_T3));
fdce N1P_1_180P_1_21P_1_I20_1_I12_1 (.q(N1P_1_NEXT_READ[11]), .d(N1P_1_180P_1_21P_1_I20_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_21P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_21P_1_I20_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_21P_1_I20_1_I13_1 (.o(N1P_1_180P_1_21P_1_I20_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_21P_1_I18_1_I8_1_I7_1 (.o(N1P_1_180P_1_21P_1_I18_1_I8_1_M0[0]), .i1(N1P_1_180P_1_21P_1_I18_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_21P_1_I18_1_I8_1_I6_1 (.o(N1P_1_180P_1_21P_1_I18_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[12]));
or2 N1P_1_180P_1_21P_1_I18_1_I8_1_I5_1 (.o(N1P_1_180P_1_21P_1_I18_1_MD[0]), .i1(N1P_1_180P_1_21P_1_I18_1_I8_1_M0[0]), .i0(N1P_1_180P_1_21P_1_I18_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_21P_1_I18_1_I9_1 (.o(N1P_1_180P_1_21P_1_I18_1_TQ[0]), .i1(N1P_1_NEXT_READ[10]), .i0(N1P_1_180P_1_21P_1_T2));
fdce N1P_1_180P_1_21P_1_I18_1_I12_1 (.q(N1P_1_NEXT_READ[10]), .d(N1P_1_180P_1_21P_1_I18_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_21P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_21P_1_I18_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_21P_1_I18_1_I13_1 (.o(N1P_1_180P_1_21P_1_I18_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and3 N1P_1_180P_1_21P_1_I21_1 (.i2(N1P_1_NEXT_READ[8]), .o(N1P_1_180P_1_21P_1_T3), .i1(N1P_1_NEXT_READ[9]), .i0(N1P_1_NEXT_READ[10]));
and4 N1P_1_180P_1_21P_1_I19_1 (.i2(N1P_1_NEXT_READ[10]), .i3(N1P_1_NEXT_READ[11]), .o(N1P_1_180P_1_UN_1_CB4CLE_21P_TC), .i1(N1P_1_NEXT_READ[9]), .i0(N1P_1_NEXT_READ[8]));
and2 N1P_1_180P_1_21P_1_I24_1 (.o(N1P_1_180P_1_21P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CLE_21P_TC), .i0(XVDD));
and2 N1P_1_180P_1_21P_1_I17_1 (.o(N1P_1_180P_1_21P_1_T2), .i1(N1P_1_NEXT_READ[8]), .i0(N1P_1_NEXT_READ[9]));
and2b1 N1P_1_180P_1_1P_1_I23_1_I8_1_I7_1 (.o(N1P_1_180P_1_1P_1_I23_1_I8_1_M0[0]), .i1(N1P_1_180P_1_1P_1_I23_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_1P_1_I23_1_I8_1_I6_1 (.o(N1P_1_180P_1_1P_1_I23_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[19]));
or2 N1P_1_180P_1_1P_1_I23_1_I8_1_I5_1 (.o(N1P_1_180P_1_1P_1_I23_1_MD[0]), .i1(N1P_1_180P_1_1P_1_I23_1_I8_1_M0[0]), .i0(N1P_1_180P_1_1P_1_I23_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_1P_1_I23_1_I9_1 (.o(N1P_1_180P_1_1P_1_I23_1_TQ[0]), .i1(N1P_1_NEXT_READ[17]), .i0(N1P_1_NEXT_READ[16]));
fdce N1P_1_180P_1_1P_1_I23_1_I12_1 (.q(N1P_1_NEXT_READ[17]), .d(N1P_1_180P_1_1P_1_I23_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_1P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_1P_1_I23_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_1P_1_I23_1_I13_1 (.o(N1P_1_180P_1_1P_1_I23_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_1P_1_I22_1_I8_1_I7_1 (.o(N1P_1_180P_1_1P_1_I22_1_I8_1_M0[0]), .i1(N1P_1_180P_1_1P_1_I22_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_1P_1_I22_1_I8_1_I6_1 (.o(N1P_1_180P_1_1P_1_I22_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[18]));
or2 N1P_1_180P_1_1P_1_I22_1_I8_1_I5_1 (.o(N1P_1_180P_1_1P_1_I22_1_MD[0]), .i1(N1P_1_180P_1_1P_1_I22_1_I8_1_M0[0]), .i0(N1P_1_180P_1_1P_1_I22_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_1P_1_I22_1_I9_1 (.o(N1P_1_180P_1_1P_1_I22_1_TQ[0]), .i1(N1P_1_NEXT_READ[16]), .i0(XVDD));
fdce N1P_1_180P_1_1P_1_I22_1_I12_1 (.q(N1P_1_NEXT_READ[16]), .d(N1P_1_180P_1_1P_1_I22_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_1P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_1P_1_I22_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_1P_1_I22_1_I13_1 (.o(N1P_1_180P_1_1P_1_I22_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_1P_1_I20_1_I8_1_I7_1 (.o(N1P_1_180P_1_1P_1_I20_1_I8_1_M0[0]), .i1(N1P_1_180P_1_1P_1_I20_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_1P_1_I20_1_I8_1_I6_1 (.o(N1P_1_180P_1_1P_1_I20_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[21]));
or2 N1P_1_180P_1_1P_1_I20_1_I8_1_I5_1 (.o(N1P_1_180P_1_1P_1_I20_1_MD[0]), .i1(N1P_1_180P_1_1P_1_I20_1_I8_1_M0[0]), .i0(N1P_1_180P_1_1P_1_I20_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_1P_1_I20_1_I9_1 (.o(N1P_1_180P_1_1P_1_I20_1_TQ[0]), .i1(N1P_1_NEXT_READ[19]), .i0(N1P_1_180P_1_1P_1_T3));
fdce N1P_1_180P_1_1P_1_I20_1_I12_1 (.q(N1P_1_NEXT_READ[19]), .d(N1P_1_180P_1_1P_1_I20_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_1P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_1P_1_I20_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_1P_1_I20_1_I13_1 (.o(N1P_1_180P_1_1P_1_I20_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_1P_1_I18_1_I8_1_I7_1 (.o(N1P_1_180P_1_1P_1_I18_1_I8_1_M0[0]), .i1(N1P_1_180P_1_1P_1_I18_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_1P_1_I18_1_I8_1_I6_1 (.o(N1P_1_180P_1_1P_1_I18_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[20]));
or2 N1P_1_180P_1_1P_1_I18_1_I8_1_I5_1 (.o(N1P_1_180P_1_1P_1_I18_1_MD[0]), .i1(N1P_1_180P_1_1P_1_I18_1_I8_1_M0[0]), .i0(N1P_1_180P_1_1P_1_I18_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_1P_1_I18_1_I9_1 (.o(N1P_1_180P_1_1P_1_I18_1_TQ[0]), .i1(N1P_1_NEXT_READ[18]), .i0(N1P_1_180P_1_1P_1_T2));
fdce N1P_1_180P_1_1P_1_I18_1_I12_1 (.q(N1P_1_NEXT_READ[18]), .d(N1P_1_180P_1_1P_1_I18_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_1P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_1P_1_I18_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_1P_1_I18_1_I13_1 (.o(N1P_1_180P_1_1P_1_I18_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and3 N1P_1_180P_1_1P_1_I21_1 (.i2(N1P_1_NEXT_READ[16]), .o(N1P_1_180P_1_1P_1_T3), .i1(N1P_1_NEXT_READ[17]), .i0(N1P_1_NEXT_READ[18]));
and4 N1P_1_180P_1_1P_1_I19_1 (.i2(N1P_1_NEXT_READ[18]), .i3(N1P_1_NEXT_READ[19]), .o(N1P_1_180P_1_1P_1_TC), .i1(N1P_1_NEXT_READ[17]), .i0(N1P_1_NEXT_READ[16]));
and2 N1P_1_180P_1_1P_1_I24_1 (.o(N1P_1_180P_1_1P_1_CEO), .i1(N1P_1_180P_1_1P_1_TC), .i0(XVDD));
and2 N1P_1_180P_1_1P_1_I17_1 (.o(N1P_1_180P_1_1P_1_T2), .i1(N1P_1_NEXT_READ[16]), .i0(N1P_1_NEXT_READ[17]));
and2b1 N1P_1_180P_1_11P_1_I23_1_I8_1_I7_1 (.o(N1P_1_180P_1_11P_1_I23_1_I8_1_M0[0]), .i1(N1P_1_180P_1_11P_1_I23_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_11P_1_I23_1_I8_1_I6_1 (.o(N1P_1_180P_1_11P_1_I23_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[15]));
or2 N1P_1_180P_1_11P_1_I23_1_I8_1_I5_1 (.o(N1P_1_180P_1_11P_1_I23_1_MD[0]), .i1(N1P_1_180P_1_11P_1_I23_1_I8_1_M0[0]), .i0(N1P_1_180P_1_11P_1_I23_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_11P_1_I23_1_I9_1 (.o(N1P_1_180P_1_11P_1_I23_1_TQ[0]), .i1(N1P_1_NEXT_READ[13]), .i0(N1P_1_NEXT_READ[12]));
fdce N1P_1_180P_1_11P_1_I23_1_I12_1 (.q(N1P_1_NEXT_READ[13]), .d(N1P_1_180P_1_11P_1_I23_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_11P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_11P_1_I23_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_11P_1_I23_1_I13_1 (.o(N1P_1_180P_1_11P_1_I23_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_11P_1_I22_1_I8_1_I7_1 (.o(N1P_1_180P_1_11P_1_I22_1_I8_1_M0[0]), .i1(N1P_1_180P_1_11P_1_I22_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_11P_1_I22_1_I8_1_I6_1 (.o(N1P_1_180P_1_11P_1_I22_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[14]));
or2 N1P_1_180P_1_11P_1_I22_1_I8_1_I5_1 (.o(N1P_1_180P_1_11P_1_I22_1_MD[0]), .i1(N1P_1_180P_1_11P_1_I22_1_I8_1_M0[0]), .i0(N1P_1_180P_1_11P_1_I22_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_11P_1_I22_1_I9_1 (.o(N1P_1_180P_1_11P_1_I22_1_TQ[0]), .i1(N1P_1_NEXT_READ[12]), .i0(XVDD));
fdce N1P_1_180P_1_11P_1_I22_1_I12_1 (.q(N1P_1_NEXT_READ[12]), .d(N1P_1_180P_1_11P_1_I22_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_11P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_11P_1_I22_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_11P_1_I22_1_I13_1 (.o(N1P_1_180P_1_11P_1_I22_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_11P_1_I20_1_I8_1_I7_1 (.o(N1P_1_180P_1_11P_1_I20_1_I8_1_M0[0]), .i1(N1P_1_180P_1_11P_1_I20_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_11P_1_I20_1_I8_1_I6_1 (.o(N1P_1_180P_1_11P_1_I20_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[17]));
or2 N1P_1_180P_1_11P_1_I20_1_I8_1_I5_1 (.o(N1P_1_180P_1_11P_1_I20_1_MD[0]), .i1(N1P_1_180P_1_11P_1_I20_1_I8_1_M0[0]), .i0(N1P_1_180P_1_11P_1_I20_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_11P_1_I20_1_I9_1 (.o(N1P_1_180P_1_11P_1_I20_1_TQ[0]), .i1(N1P_1_NEXT_READ[15]), .i0(N1P_1_180P_1_11P_1_T3));
fdce N1P_1_180P_1_11P_1_I20_1_I12_1 (.q(N1P_1_NEXT_READ[15]), .d(N1P_1_180P_1_11P_1_I20_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_11P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_11P_1_I20_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_11P_1_I20_1_I13_1 (.o(N1P_1_180P_1_11P_1_I20_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and2b1 N1P_1_180P_1_11P_1_I18_1_I8_1_I7_1 (.o(N1P_1_180P_1_11P_1_I18_1_I8_1_M0[0]), .i1(N1P_1_180P_1_11P_1_I18_1_TQ[0]), .i0(N1P_1_SEL1));
and2 N1P_1_180P_1_11P_1_I18_1_I8_1_I6_1 (.o(N1P_1_180P_1_11P_1_I18_1_I8_1_M1[0]), .i1(N1P_1_SEL1), .i0(BBA[16]));
or2 N1P_1_180P_1_11P_1_I18_1_I8_1_I5_1 (.o(N1P_1_180P_1_11P_1_I18_1_MD[0]), .i1(N1P_1_180P_1_11P_1_I18_1_I8_1_M0[0]), .i0(N1P_1_180P_1_11P_1_I18_1_I8_1_M1[0]));
xor2 N1P_1_180P_1_11P_1_I18_1_I9_1 (.o(N1P_1_180P_1_11P_1_I18_1_TQ[0]), .i1(N1P_1_NEXT_READ[14]), .i0(N1P_1_180P_1_11P_1_T2));
fdce N1P_1_180P_1_11P_1_I18_1_I12_1 (.q(N1P_1_NEXT_READ[14]), .d(N1P_1_180P_1_11P_1_I18_1_MD[0]), .c(N1P_1_180P_1_UN_1_CB4CLE_11P_C), .clr(N1P_1_FIFO_RESET), .ce(N1P_1_180P_1_11P_1_I18_1_L_CE), .gr(RESET_n));
or2 N1P_1_180P_1_11P_1_I18_1_I13_1 (.o(N1P_1_180P_1_11P_1_I18_1_L_CE), .i1(N1P_1_SEL1), .i0(XVDD));
and3 N1P_1_180P_1_11P_1_I21_1 (.i2(N1P_1_NEXT_READ[12]), .o(N1P_1_180P_1_11P_1_T3), .i1(N1P_1_NEXT_READ[13]), .i0(N1P_1_NEXT_READ[14]));
and4 N1P_1_180P_1_11P_1_I19_1 (.i2(N1P_1_NEXT_READ[14]), .i3(N1P_1_NEXT_READ[15]), .o(N1P_1_180P_1_UN_1_CB4CLE_11P_TC), .i1(N1P_1_NEXT_READ[13]), .i0(N1P_1_NEXT_READ[12]));
and2 N1P_1_180P_1_11P_1_I24_1 (.o(N1P_1_180P_1_11P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CLE_11P_TC), .i0(XVDD));
and2 N1P_1_180P_1_11P_1_I17_1 (.o(N1P_1_180P_1_11P_1_T2), .i1(N1P_1_NEXT_READ[12]), .i0(N1P_1_NEXT_READ[13]));
xor2 N1P_1_180P_1_71P_1_I19_1_I8_1 (.o(N1P_1_180P_1_71P_1_I19_1_TQ[0]), .i1(BWR_ADD[16]), .i0(N1P_1_180P_1_71P_1_T2));
fdce N1P_1_180P_1_71P_1_I19_1_I7_1 (.q(BWR_ADD[16]), .d(N1P_1_180P_1_71P_1_I19_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_71P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_71P_1_I18_1_I8_1 (.o(N1P_1_180P_1_71P_1_I18_1_TQ[0]), .i1(BWR_ADD[15]), .i0(BWR_ADD[14]));
fdce N1P_1_180P_1_71P_1_I18_1_I7_1 (.q(BWR_ADD[15]), .d(N1P_1_180P_1_71P_1_I18_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_71P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_71P_1_I12_1_I8_1 (.o(N1P_1_180P_1_71P_1_I12_1_TQ[0]), .i1(BWR_ADD[14]), .i0(XVDD));
fdce N1P_1_180P_1_71P_1_I12_1_I7_1 (.q(BWR_ADD[14]), .d(N1P_1_180P_1_71P_1_I12_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_71P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_71P_1_I11_1_I8_1 (.o(N1P_1_180P_1_71P_1_I11_1_TQ[0]), .i1(BWR_ADD[17]), .i0(N1P_1_180P_1_71P_1_T3));
fdce N1P_1_180P_1_71P_1_I11_1_I7_1 (.q(BWR_ADD[17]), .d(N1P_1_180P_1_71P_1_I11_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_71P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
and3 N1P_1_180P_1_71P_1_I13_1 (.i2(BWR_ADD[14]), .o(N1P_1_180P_1_71P_1_T3), .i1(BWR_ADD[15]), .i0(BWR_ADD[16]));
and4 N1P_1_180P_1_71P_1_I10_1 (.i2(BWR_ADD[15]), .i3(BWR_ADD[14]), .o(N1P_1_180P_1_UN_1_CB4CE_71P_TC), .i1(BWR_ADD[16]), .i0(BWR_ADD[17]));
and2 N1P_1_180P_1_71P_1_I16_1 (.o(N1P_1_180P_1_71P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CE_71P_TC), .i0(XVDD));
and2 N1P_1_180P_1_71P_1_I14_1 (.o(N1P_1_180P_1_71P_1_T2), .i1(BWR_ADD[14]), .i0(BWR_ADD[15]));
xor2 N1P_1_180P_1_77P_1_I19_1_I8_1 (.o(N1P_1_180P_1_77P_1_I19_1_TQ[0]), .i1(BWR_ADD[20]), .i0(N1P_1_180P_1_77P_1_T2));
fdce N1P_1_180P_1_77P_1_I19_1_I7_1 (.q(BWR_ADD[20]), .d(N1P_1_180P_1_77P_1_I19_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_77P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_77P_1_I18_1_I8_1 (.o(N1P_1_180P_1_77P_1_I18_1_TQ[0]), .i1(BWR_ADD[19]), .i0(BWR_ADD[18]));
fdce N1P_1_180P_1_77P_1_I18_1_I7_1 (.q(BWR_ADD[19]), .d(N1P_1_180P_1_77P_1_I18_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_77P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_77P_1_I12_1_I8_1 (.o(N1P_1_180P_1_77P_1_I12_1_TQ[0]), .i1(BWR_ADD[18]), .i0(XVDD));
fdce N1P_1_180P_1_77P_1_I12_1_I7_1 (.q(BWR_ADD[18]), .d(N1P_1_180P_1_77P_1_I12_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_77P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_77P_1_I11_1_I8_1 (.o(N1P_1_180P_1_77P_1_I11_1_TQ[0]), .i1(BWR_ADD[21]), .i0(N1P_1_180P_1_77P_1_T3));
fdce N1P_1_180P_1_77P_1_I11_1_I7_1 (.q(BWR_ADD[21]), .d(N1P_1_180P_1_77P_1_I11_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_77P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
and3 N1P_1_180P_1_77P_1_I13_1 (.i2(BWR_ADD[18]), .o(N1P_1_180P_1_77P_1_T3), .i1(BWR_ADD[19]), .i0(BWR_ADD[20]));
and4 N1P_1_180P_1_77P_1_I10_1 (.i2(BWR_ADD[19]), .i3(BWR_ADD[18]), .o(N1P_1_180P_1_77P_1_TC), .i1(BWR_ADD[20]), .i0(BWR_ADD[21]));
and2 N1P_1_180P_1_77P_1_I16_1 (.o(N1P_1_180P_1_77P_1_CEO), .i1(N1P_1_180P_1_77P_1_TC), .i0(XVDD));
and2 N1P_1_180P_1_77P_1_I14_1 (.o(N1P_1_180P_1_77P_1_T2), .i1(BWR_ADD[18]), .i0(BWR_ADD[19]));
xor2 N1P_1_180P_1_65P_1_I19_1_I8_1 (.o(N1P_1_180P_1_65P_1_I19_1_TQ[0]), .i1(BWR_ADD[12]), .i0(N1P_1_180P_1_65P_1_T2));
fdce N1P_1_180P_1_65P_1_I19_1_I7_1 (.q(BWR_ADD[12]), .d(N1P_1_180P_1_65P_1_I19_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_65P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_65P_1_I18_1_I8_1 (.o(N1P_1_180P_1_65P_1_I18_1_TQ[0]), .i1(BWR_ADD[11]), .i0(BWR_ADD[10]));
fdce N1P_1_180P_1_65P_1_I18_1_I7_1 (.q(BWR_ADD[11]), .d(N1P_1_180P_1_65P_1_I18_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_65P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_65P_1_I12_1_I8_1 (.o(N1P_1_180P_1_65P_1_I12_1_TQ[0]), .i1(BWR_ADD[10]), .i0(XVDD));
fdce N1P_1_180P_1_65P_1_I12_1_I7_1 (.q(BWR_ADD[10]), .d(N1P_1_180P_1_65P_1_I12_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_65P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_65P_1_I11_1_I8_1 (.o(N1P_1_180P_1_65P_1_I11_1_TQ[0]), .i1(BWR_ADD[13]), .i0(N1P_1_180P_1_65P_1_T3));
fdce N1P_1_180P_1_65P_1_I11_1_I7_1 (.q(BWR_ADD[13]), .d(N1P_1_180P_1_65P_1_I11_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_65P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
and3 N1P_1_180P_1_65P_1_I13_1 (.i2(BWR_ADD[10]), .o(N1P_1_180P_1_65P_1_T3), .i1(BWR_ADD[11]), .i0(BWR_ADD[12]));
and4 N1P_1_180P_1_65P_1_I10_1 (.i2(BWR_ADD[11]), .i3(BWR_ADD[10]), .o(N1P_1_180P_1_UN_1_CB4CE_65P_TC), .i1(BWR_ADD[12]), .i0(BWR_ADD[13]));
and2 N1P_1_180P_1_65P_1_I16_1 (.o(N1P_1_180P_1_65P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CE_65P_TC), .i0(XVDD));
and2 N1P_1_180P_1_65P_1_I14_1 (.o(N1P_1_180P_1_65P_1_T2), .i1(BWR_ADD[10]), .i0(BWR_ADD[11]));
xor2 N1P_1_180P_1_59P_1_I19_1_I8_1 (.o(N1P_1_180P_1_59P_1_I19_1_TQ[0]), .i1(BWR_ADD[8]), .i0(N1P_1_180P_1_59P_1_T2));
fdce N1P_1_180P_1_59P_1_I19_1_I7_1 (.q(BWR_ADD[8]), .d(N1P_1_180P_1_59P_1_I19_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_59P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_59P_1_I18_1_I8_1 (.o(N1P_1_180P_1_59P_1_I18_1_TQ[0]), .i1(BWR_ADD[7]), .i0(BWR_ADD[6]));
fdce N1P_1_180P_1_59P_1_I18_1_I7_1 (.q(BWR_ADD[7]), .d(N1P_1_180P_1_59P_1_I18_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_59P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_59P_1_I12_1_I8_1 (.o(N1P_1_180P_1_59P_1_I12_1_TQ[0]), .i1(BWR_ADD[6]), .i0(XVDD));
fdce N1P_1_180P_1_59P_1_I12_1_I7_1 (.q(BWR_ADD[6]), .d(N1P_1_180P_1_59P_1_I12_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_59P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_59P_1_I11_1_I8_1 (.o(N1P_1_180P_1_59P_1_I11_1_TQ[0]), .i1(BWR_ADD[9]), .i0(N1P_1_180P_1_59P_1_T3));
fdce N1P_1_180P_1_59P_1_I11_1_I7_1 (.q(BWR_ADD[9]), .d(N1P_1_180P_1_59P_1_I11_1_TQ[0]), .c(N1P_1_180P_1_UN_1_CB4CE_59P_C), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
and3 N1P_1_180P_1_59P_1_I13_1 (.i2(BWR_ADD[6]), .o(N1P_1_180P_1_59P_1_T3), .i1(BWR_ADD[7]), .i0(BWR_ADD[8]));
and4 N1P_1_180P_1_59P_1_I10_1 (.i2(BWR_ADD[7]), .i3(BWR_ADD[6]), .o(N1P_1_180P_1_UN_1_CB4CE_59P_TC), .i1(BWR_ADD[8]), .i0(BWR_ADD[9]));
and2 N1P_1_180P_1_59P_1_I16_1 (.o(N1P_1_180P_1_59P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CE_59P_TC), .i0(XVDD));
and2 N1P_1_180P_1_59P_1_I14_1 (.o(N1P_1_180P_1_59P_1_T2), .i1(BWR_ADD[6]), .i0(BWR_ADD[7]));
xor2 N1P_1_180P_1_53P_1_I19_1_I8_1 (.o(N1P_1_180P_1_53P_1_I19_1_TQ[0]), .i1(BWR_ADD[4]), .i0(N1P_1_180P_1_53P_1_T2));
fdce N1P_1_180P_1_53P_1_I19_1_I7_1 (.q(BWR_ADD[4]), .d(N1P_1_180P_1_53P_1_I19_1_TQ[0]), .c(MEMACK2_n), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_53P_1_I18_1_I8_1 (.o(N1P_1_180P_1_53P_1_I18_1_TQ[0]), .i1(BWR_ADD[3]), .i0(BWR_ADD[2]));
fdce N1P_1_180P_1_53P_1_I18_1_I7_1 (.q(BWR_ADD[3]), .d(N1P_1_180P_1_53P_1_I18_1_TQ[0]), .c(MEMACK2_n), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_53P_1_I12_1_I8_1 (.o(N1P_1_180P_1_53P_1_I12_1_TQ[0]), .i1(BWR_ADD[2]), .i0(XVDD));
fdce N1P_1_180P_1_53P_1_I12_1_I7_1 (.q(BWR_ADD[2]), .d(N1P_1_180P_1_53P_1_I12_1_TQ[0]), .c(MEMACK2_n), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
xor2 N1P_1_180P_1_53P_1_I11_1_I8_1 (.o(N1P_1_180P_1_53P_1_I11_1_TQ[0]), .i1(BWR_ADD[5]), .i0(N1P_1_180P_1_53P_1_T3));
fdce N1P_1_180P_1_53P_1_I11_1_I7_1 (.q(BWR_ADD[5]), .d(N1P_1_180P_1_53P_1_I11_1_TQ[0]), .c(MEMACK2_n), .clr(N1P_1_FIFO_RESET), .ce(XVDD), .gr(RESET_n));
and3 N1P_1_180P_1_53P_1_I13_1 (.i2(BWR_ADD[2]), .o(N1P_1_180P_1_53P_1_T3), .i1(BWR_ADD[3]), .i0(BWR_ADD[4]));
and4 N1P_1_180P_1_53P_1_I10_1 (.i2(BWR_ADD[3]), .i3(BWR_ADD[2]), .o(N1P_1_180P_1_UN_1_CB4CE_53P_TC), .i1(BWR_ADD[4]), .i0(BWR_ADD[5]));
and2 N1P_1_180P_1_53P_1_I16_1 (.o(N1P_1_180P_1_53P_1_CEO), .i1(N1P_1_180P_1_UN_1_CB4CE_53P_TC), .i0(XVDD));
and2 N1P_1_180P_1_53P_1_I14_1 (.o(N1P_1_180P_1_53P_1_T2), .i1(BWR_ADD[2]), .i0(BWR_ADD[3]));
inv N1P_1_180P_1_64P_1 (.i(N1P_1_180P_1_UN_1_CB4CE_59P_TC), .o(N1P_1_180P_1_UN_1_CB4CE_65P_C));
inv N1P_1_180P_1_70P_1 (.i(N1P_1_180P_1_UN_1_CB4CE_65P_TC), .o(N1P_1_180P_1_UN_1_CB4CE_71P_C));
inv N1P_1_180P_1_76P_1 (.i(N1P_1_180P_1_UN_1_CB4CE_71P_TC), .o(N1P_1_180P_1_UN_1_CB4CE_77P_C));
inv N1P_1_180P_1_58P_1 (.i(N1P_1_180P_1_UN_1_CB4CE_53P_TC), .o(N1P_1_180P_1_UN_1_CB4CE_59P_C));
inv N1P_1_180P_1_40P_1 (.i(N1P_1_180P_1_UN_1_CB4CLE_41P_TC), .o(N1P_1_180P_1_UN_1_CB4CLE_31P_C));
inv N1P_1_180P_1_30P_1 (.i(N1P_1_180P_1_UN_1_CB4CLE_31P_TC), .o(N1P_1_180P_1_UN_1_CB4CLE_21P_C));
inv N1P_1_180P_1_20P_1 (.i(N1P_1_180P_1_UN_1_CB4CLE_21P_TC), .o(N1P_1_180P_1_UN_1_CB4CLE_11P_C));
inv N1P_1_180P_1_10P_1 (.i(N1P_1_180P_1_UN_1_CB4CLE_11P_TC), .o(N1P_1_180P_1_UN_1_CB4CLE_1P_C));
xnor2 N1P_1_179P_1_70P_1_I15_1 (.o(N1P_1_179P_1_70P_1_AB1[0]), .i1(N1P_1_NEXT_READ[13]), .i0(BWR_ADD[15]));
xnor2 N1P_1_179P_1_70P_1_I14_1 (.o(N1P_1_179P_1_70P_1_AB0[0]), .i1(N1P_1_NEXT_READ[12]), .i0(BWR_ADD[14]));
xnor2 N1P_1_179P_1_70P_1_I12_1 (.o(N1P_1_179P_1_70P_1_AB2[0]), .i1(N1P_1_NEXT_READ[14]), .i0(BWR_ADD[16]));
xnor2 N1P_1_179P_1_70P_1_I11_1 (.o(N1P_1_179P_1_70P_1_AB3[0]), .i1(N1P_1_NEXT_READ[15]), .i0(BWR_ADD[17]));
and4 N1P_1_179P_1_70P_1_I10_1 (.i2(N1P_1_179P_1_70P_1_AB1[0]), .i3(N1P_1_179P_1_70P_1_AB0[0]), .o(N1P_1_179P_1_UN_1_AND5_2P_I3), .i1(N1P_1_179P_1_70P_1_AB2[0]), .i0(N1P_1_179P_1_70P_1_AB3[0]));
xnor2 N1P_1_179P_1_62P_1_I15_1 (.o(N1P_1_179P_1_62P_1_AB1[0]), .i1(N1P_1_NEXT_READ[5]), .i0(BWR_ADD[7]));
xnor2 N1P_1_179P_1_62P_1_I14_1 (.o(N1P_1_179P_1_62P_1_AB0[0]), .i1(N1P_1_NEXT_READ[4]), .i0(BWR_ADD[6]));
xnor2 N1P_1_179P_1_62P_1_I12_1 (.o(N1P_1_179P_1_62P_1_AB2[0]), .i1(N1P_1_NEXT_READ[6]), .i0(BWR_ADD[8]));
xnor2 N1P_1_179P_1_62P_1_I11_1 (.o(N1P_1_179P_1_62P_1_AB3[0]), .i1(N1P_1_NEXT_READ[7]), .i0(BWR_ADD[9]));
and4 N1P_1_179P_1_62P_1_I10_1 (.i2(N1P_1_179P_1_62P_1_AB1[0]), .i3(N1P_1_179P_1_62P_1_AB0[0]), .o(N1P_1_179P_1_UN_1_AND5_2P_I1), .i1(N1P_1_179P_1_62P_1_AB2[0]), .i0(N1P_1_179P_1_62P_1_AB3[0]));
xnor2 N1P_1_179P_1_74P_1_I15_1 (.o(N1P_1_179P_1_74P_1_AB1[0]), .i1(N1P_1_NEXT_READ[17]), .i0(BWR_ADD[19]));
xnor2 N1P_1_179P_1_74P_1_I14_1 (.o(N1P_1_179P_1_74P_1_AB0[0]), .i1(N1P_1_NEXT_READ[16]), .i0(BWR_ADD[18]));
xnor2 N1P_1_179P_1_74P_1_I12_1 (.o(N1P_1_179P_1_74P_1_AB2[0]), .i1(N1P_1_NEXT_READ[18]), .i0(BWR_ADD[20]));
xnor2 N1P_1_179P_1_74P_1_I11_1 (.o(N1P_1_179P_1_74P_1_AB3[0]), .i1(N1P_1_NEXT_READ[19]), .i0(BWR_ADD[21]));
and4 N1P_1_179P_1_74P_1_I10_1 (.i2(N1P_1_179P_1_74P_1_AB1[0]), .i3(N1P_1_179P_1_74P_1_AB0[0]), .o(N1P_1_179P_1_UN_1_AND5_2P_I4), .i1(N1P_1_179P_1_74P_1_AB2[0]), .i0(N1P_1_179P_1_74P_1_AB3[0]));
xnor2 N1P_1_179P_1_66P_1_I15_1 (.o(N1P_1_179P_1_66P_1_AB1[0]), .i1(N1P_1_NEXT_READ[9]), .i0(BWR_ADD[11]));
xnor2 N1P_1_179P_1_66P_1_I14_1 (.o(N1P_1_179P_1_66P_1_AB0[0]), .i1(N1P_1_NEXT_READ[8]), .i0(BWR_ADD[10]));
xnor2 N1P_1_179P_1_66P_1_I12_1 (.o(N1P_1_179P_1_66P_1_AB2[0]), .i1(N1P_1_NEXT_READ[10]), .i0(BWR_ADD[12]));
xnor2 N1P_1_179P_1_66P_1_I11_1 (.o(N1P_1_179P_1_66P_1_AB3[0]), .i1(N1P_1_NEXT_READ[11]), .i0(BWR_ADD[13]));
and4 N1P_1_179P_1_66P_1_I10_1 (.i2(N1P_1_179P_1_66P_1_AB1[0]), .i3(N1P_1_179P_1_66P_1_AB0[0]), .o(N1P_1_179P_1_UN_1_AND5_2P_I2), .i1(N1P_1_179P_1_66P_1_AB2[0]), .i0(N1P_1_179P_1_66P_1_AB3[0]));
xnor2 N1P_1_179P_1_58P_1_I15_1 (.o(N1P_1_179P_1_58P_1_AB1[0]), .i1(N1P_1_NEXT_READ[1]), .i0(BWR_ADD[3]));
xnor2 N1P_1_179P_1_58P_1_I14_1 (.o(N1P_1_179P_1_58P_1_AB0[0]), .i1(N1P_1_NEXT_READ[0]), .i0(BWR_ADD[2]));
xnor2 N1P_1_179P_1_58P_1_I12_1 (.o(N1P_1_179P_1_58P_1_AB2[0]), .i1(N1P_1_NEXT_READ[2]), .i0(BWR_ADD[4]));
xnor2 N1P_1_179P_1_58P_1_I11_1 (.o(N1P_1_179P_1_58P_1_AB3[0]), .i1(N1P_1_NEXT_READ[3]), .i0(BWR_ADD[5]));
and4 N1P_1_179P_1_58P_1_I10_1 (.i2(N1P_1_179P_1_58P_1_AB1[0]), .i3(N1P_1_179P_1_58P_1_AB0[0]), .o(N1P_1_179P_1_UN_1_AND5_2P_I0), .i1(N1P_1_179P_1_58P_1_AB2[0]), .i0(N1P_1_179P_1_58P_1_AB3[0]));
or5 N1P_1_179P_1_47P_1_I32_1 (.i2(N1P_1_179P_1_47P_1_AB3), .i3(N1P_1_179P_1_47P_1_AB1), .i4(N1P_1_179P_1_47P_1_AG_7), .o(N1P_1_179P_1_UN_1_X74_L85_39P_ALBI), .i1(N1P_1_179P_1_47P_1_AB5), .i0(N1P_1_179P_1_47P_1_AB7));
or5 N1P_1_179P_1_47P_1_I24_1 (.i2(N1P_1_179P_1_47P_1_AB2), .i3(N1P_1_179P_1_47P_1_AB0), .i4(N1P_1_179P_1_47P_1_AL_7), .o(N1P_1_179P_1_UN_1_X74_L85_39P_AGBI), .i1(N1P_1_179P_1_47P_1_AB4), .i0(N1P_1_179P_1_47P_1_AB6));
and2b1 N1P_1_179P_1_47P_1_I41_1 (.o(N1P_1_179P_1_47P_1_A_B0), .i1(N1P_1_LAST_WRITE[0]), .i0(N1P_1_LAST_READ[0]));
and2b1 N1P_1_179P_1_47P_1_I40_1 (.o(N1P_1_179P_1_47P_1_A_B5), .i1(N1P_1_LAST_READ[2]), .i0(N1P_1_LAST_WRITE[2]));
and2b1 N1P_1_179P_1_47P_1_I38_1 (.o(N1P_1_179P_1_47P_1_A_B2), .i1(N1P_1_LAST_WRITE[1]), .i0(N1P_1_LAST_READ[1]));
and2b1 N1P_1_179P_1_47P_1_I37_1 (.o(N1P_1_179P_1_47P_1_A_B7), .i1(N1P_1_LAST_READ[3]), .i0(N1P_1_LAST_WRITE[3]));
and2b1 N1P_1_179P_1_47P_1_I36_1 (.o(N1P_1_179P_1_47P_1_AB6), .i1(N1P_1_LAST_READ[3]), .i0(N1P_1_LAST_WRITE[3]));
and2b1 N1P_1_179P_1_47P_1_I30_1 (.o(N1P_1_179P_1_47P_1_AB7), .i1(N1P_1_LAST_WRITE[3]), .i0(N1P_1_LAST_READ[3]));
and2b1 N1P_1_179P_1_47P_1_I29_1 (.o(N1P_1_179P_1_47P_1_A_B1), .i1(N1P_1_LAST_READ[0]), .i0(N1P_1_LAST_WRITE[0]));
and2b1 N1P_1_179P_1_47P_1_I28_1 (.o(N1P_1_179P_1_47P_1_A_B4), .i1(N1P_1_LAST_WRITE[2]), .i0(N1P_1_LAST_READ[2]));
and2b1 N1P_1_179P_1_47P_1_I26_1 (.o(N1P_1_179P_1_47P_1_A_B6), .i1(N1P_1_LAST_WRITE[3]), .i0(N1P_1_LAST_READ[3]));
and2b1 N1P_1_179P_1_47P_1_I22_1 (.o(N1P_1_179P_1_47P_1_A_B3), .i1(N1P_1_LAST_READ[1]), .i0(N1P_1_LAST_WRITE[1]));
and4b1 N1P_1_179P_1_47P_1_I21_1 (.i3(N1P_1_179P_1_47P_1_NA_B5), .i2(N1P_1_LAST_WRITE[1]), .o(N1P_1_179P_1_47P_1_AB3), .i1(N1P_1_179P_1_47P_1_NA_B7), .i0(N1P_1_LAST_READ[1]));
and4b1 N1P_1_179P_1_47P_1_I20_1 (.i3(N1P_1_179P_1_47P_1_NA_B5), .i2(N1P_1_LAST_READ[1]), .o(N1P_1_179P_1_47P_1_AB2), .i1(N1P_1_179P_1_47P_1_NA_B7), .i0(N1P_1_LAST_WRITE[1]));
and5b1 N1P_1_179P_1_47P_1_I25_1 (.i4(N1P_1_179P_1_47P_1_NA_B5), .i3(N1P_1_179P_1_47P_1_NA_B3), .i2(N1P_1_LAST_READ[0]), .o(N1P_1_179P_1_47P_1_AB0), .i1(N1P_1_179P_1_47P_1_NA_B7), .i0(N1P_1_LAST_WRITE[0]));
and5b1 N1P_1_179P_1_47P_1_I16_1 (.i4(N1P_1_179P_1_47P_1_NA_B5), .i3(N1P_1_179P_1_47P_1_NA_B3), .i2(N1P_1_LAST_WRITE[0]), .o(N1P_1_179P_1_47P_1_AB1), .i1(N1P_1_179P_1_47P_1_NA_B7), .i0(N1P_1_LAST_READ[0]));
and3b1 N1P_1_179P_1_47P_1_I27_1 (.i2(N1P_1_LAST_READ[2]), .o(N1P_1_179P_1_47P_1_AB4), .i1(N1P_1_179P_1_47P_1_NA_B7), .i0(N1P_1_LAST_WRITE[2]));
and3b1 N1P_1_179P_1_47P_1_I15_1 (.i2(N1P_1_LAST_WRITE[2]), .o(N1P_1_179P_1_47P_1_AB5), .i1(N1P_1_179P_1_47P_1_NA_B7), .i0(N1P_1_LAST_READ[2]));
and5 N1P_1_179P_1_47P_1_I23_1 (.i2(N1P_1_179P_1_47P_1_NA_B3), .i3(N1P_1_179P_1_47P_1_NA_B1), .i4(XVDD), .o(N1P_1_179P_1_UN_1_X74_L85_39P_AEBI), .i1(N1P_1_179P_1_47P_1_NA_B5), .i0(N1P_1_179P_1_47P_1_NA_B7));
and5 N1P_1_179P_1_47P_1_I19_1 (.i2(N1P_1_179P_1_47P_1_NA_B3), .i3(N1P_1_179P_1_47P_1_NA_B1), .i4(XGND), .o(N1P_1_179P_1_47P_1_AL_7), .i1(N1P_1_179P_1_47P_1_NA_B5), .i0(N1P_1_179P_1_47P_1_NA_B7));
and5 N1P_1_179P_1_47P_1_I18_1 (.i2(N1P_1_179P_1_47P_1_NA_B3), .i3(N1P_1_179P_1_47P_1_NA_B1), .i4(XGND), .o(N1P_1_179P_1_47P_1_AG_7), .i1(N1P_1_179P_1_47P_1_NA_B5), .i0(N1P_1_179P_1_47P_1_NA_B7));
nor2 N1P_1_179P_1_47P_1_I39_1 (.o(N1P_1_179P_1_47P_1_NA_B3), .i1(N1P_1_179P_1_47P_1_A_B2), .i0(N1P_1_179P_1_47P_1_A_B3));
nor2 N1P_1_179P_1_47P_1_I35_1 (.o(N1P_1_179P_1_47P_1_NA_B1), .i1(N1P_1_179P_1_47P_1_A_B0), .i0(N1P_1_179P_1_47P_1_A_B1));
nor2 N1P_1_179P_1_47P_1_I31_1 (.o(N1P_1_179P_1_47P_1_NA_B7), .i1(N1P_1_179P_1_47P_1_A_B6), .i0(N1P_1_179P_1_47P_1_A_B7));
nor2 N1P_1_179P_1_47P_1_I17_1 (.o(N1P_1_179P_1_47P_1_NA_B5), .i1(N1P_1_179P_1_47P_1_A_B4), .i0(N1P_1_179P_1_47P_1_A_B5));
or5 N1P_1_179P_1_39P_1_I32_1 (.i2(N1P_1_179P_1_39P_1_AB3), .i3(N1P_1_179P_1_39P_1_AB1), .i4(N1P_1_179P_1_39P_1_AG_7), .o(N1P_1_179P_1_UN_1_AND2_41P_I0), .i1(N1P_1_179P_1_39P_1_AB5), .i0(N1P_1_179P_1_39P_1_AB7));
or5 N1P_1_179P_1_39P_1_I24_1 (.i2(N1P_1_179P_1_39P_1_AB2), .i3(N1P_1_179P_1_39P_1_AB0), .i4(N1P_1_179P_1_39P_1_AL_7), .o(N1P_1_179P_1_UN_1_OR2_40P_I1), .i1(N1P_1_179P_1_39P_1_AB4), .i0(N1P_1_179P_1_39P_1_AB6));
and2b1 N1P_1_179P_1_39P_1_I41_1 (.o(N1P_1_179P_1_39P_1_A_B0), .i1(N1P_1_179P_1_UN_1_X74_L85_39P_B0), .i0(N1P_1_179P_1_UN_1_X74_L85_39P_A0));
and2b1 N1P_1_179P_1_39P_1_I40_1 (.o(N1P_1_179P_1_39P_1_A_B5), .i1(N1P_1_179P_1_UN_1_X74_L85_26P_AGBO), .i0(N1P_1_179P_1_UN_1_X74_L85_26P_ALBO));
and2b1 N1P_1_179P_1_39P_1_I38_1 (.o(N1P_1_179P_1_39P_1_A_B2), .i1(N1P_1_179P_1_UN_1_X74_L85_15P_ALBO), .i0(N1P_1_179P_1_UN_1_X74_L85_15P_AGBO));
and2b1 N1P_1_179P_1_39P_1_I37_1 (.o(N1P_1_179P_1_39P_1_A_B7), .i1(N1P_1_179P_1_UN_1_X74_L85_37P_AGBO), .i0(N1P_1_179P_1_UN_1_X74_L85_37P_ALBO));
and2b1 N1P_1_179P_1_39P_1_I36_1 (.o(N1P_1_179P_1_39P_1_AB6), .i1(N1P_1_179P_1_UN_1_X74_L85_37P_AGBO), .i0(N1P_1_179P_1_UN_1_X74_L85_37P_ALBO));
and2b1 N1P_1_179P_1_39P_1_I30_1 (.o(N1P_1_179P_1_39P_1_AB7), .i1(N1P_1_179P_1_UN_1_X74_L85_37P_ALBO), .i0(N1P_1_179P_1_UN_1_X74_L85_37P_AGBO));
and2b1 N1P_1_179P_1_39P_1_I29_1 (.o(N1P_1_179P_1_39P_1_A_B1), .i1(N1P_1_179P_1_UN_1_X74_L85_39P_A0), .i0(N1P_1_179P_1_UN_1_X74_L85_39P_B0));
and2b1 N1P_1_179P_1_39P_1_I28_1 (.o(N1P_1_179P_1_39P_1_A_B4), .i1(N1P_1_179P_1_UN_1_X74_L85_26P_ALBO), .i0(N1P_1_179P_1_UN_1_X74_L85_26P_AGBO));
and2b1 N1P_1_179P_1_39P_1_I26_1 (.o(N1P_1_179P_1_39P_1_A_B6), .i1(N1P_1_179P_1_UN_1_X74_L85_37P_ALBO), .i0(N1P_1_179P_1_UN_1_X74_L85_37P_AGBO));
and2b1 N1P_1_179P_1_39P_1_I22_1 (.o(N1P_1_179P_1_39P_1_A_B3), .i1(N1P_1_179P_1_UN_1_X74_L85_15P_AGBO), .i0(N1P_1_179P_1_UN_1_X74_L85_15P_ALBO));
and4b1 N1P_1_179P_1_39P_1_I21_1 (.i3(N1P_1_179P_1_39P_1_NA_B5), .i2(N1P_1_179P_1_UN_1_X74_L85_15P_ALBO), .o(N1P_1_179P_1_39P_1_AB3), .i1(N1P_1_179P_1_39P_1_NA_B7), .i0(N1P_1_179P_1_UN_1_X74_L85_15P_AGBO));
and4b1 N1P_1_179P_1_39P_1_I20_1 (.i3(N1P_1_179P_1_39P_1_NA_B5), .i2(N1P_1_179P_1_UN_1_X74_L85_15P_AGBO), .o(N1P_1_179P_1_39P_1_AB2), .i1(N1P_1_179P_1_39P_1_NA_B7), .i0(N1P_1_179P_1_UN_1_X74_L85_15P_ALBO));
and5b1 N1P_1_179P_1_39P_1_I25_1 (.i4(N1P_1_179P_1_39P_1_NA_B5), .i3(N1P_1_179P_1_39P_1_NA_B3), .i2(N1P_1_179P_1_UN_1_X74_L85_39P_A0), .o(N1P_1_179P_1_39P_1_AB0), .i1(N1P_1_179P_1_39P_1_NA_B7), .i0(N1P_1_179P_1_UN_1_X74_L85_39P_B0));
and5b1 N1P_1_179P_1_39P_1_I16_1 (.i4(N1P_1_179P_1_39P_1_NA_B5), .i3(N1P_1_179P_1_39P_1_NA_B3), .i2(N1P_1_179P_1_UN_1_X74_L85_39P_B0), .o(N1P_1_179P_1_39P_1_AB1), .i1(N1P_1_179P_1_39P_1_NA_B7), .i0(N1P_1_179P_1_UN_1_X74_L85_39P_A0));
and3b1 N1P_1_179P_1_39P_1_I27_1 (.i2(N1P_1_179P_1_UN_1_X74_L85_26P_AGBO), .o(N1P_1_179P_1_39P_1_AB4), .i1(N1P_1_179P_1_39P_1_NA_B7), .i0(N1P_1_179P_1_UN_1_X74_L85_26P_ALBO));
and3b1 N1P_1_179P_1_39P_1_I15_1 (.i2(N1P_1_179P_1_UN_1_X74_L85_26P_ALBO), .o(N1P_1_179P_1_39P_1_AB5), .i1(N1P_1_179P_1_39P_1_NA_B7), .i0(N1P_1_179P_1_UN_1_X74_L85_26P_AGBO));
and5 N1P_1_179P_1_39P_1_I23_1 (.i2(N1P_1_179P_1_39P_1_NA_B3), .i3(N1P_1_179P_1_39P_1_NA_B1), .i4(N1P_1_179P_1_UN_1_X74_L85_39P_AEBI), .o(N1P_1_179P_1_UN_1_OR2_40P_I0), .i1(N1P_1_179P_1_39P_1_NA_B5), .i0(N1P_1_179P_1_39P_1_NA_B7));
and5 N1P_1_179P_1_39P_1_I19_1 (.i2(N1P_1_179P_1_39P_1_NA_B3), .i3(N1P_1_179P_1_39P_1_NA_B1), .i4(N1P_1_179P_1_UN_1_X74_L85_39P_AGBI), .o(N1P_1_179P_1_39P_1_AL_7), .i1(N1P_1_179P_1_39P_1_NA_B5), .i0(N1P_1_179P_1_39P_1_NA_B7));
and5 N1P_1_179P_1_39P_1_I18_1 (.i2(N1P_1_179P_1_39P_1_NA_B3), .i3(N1P_1_179P_1_39P_1_NA_B1), .i4(N1P_1_179P_1_UN_1_X74_L85_39P_ALBI), .o(N1P_1_179P_1_39P_1_AG_7), .i1(N1P_1_179P_1_39P_1_NA_B5), .i0(N1P_1_179P_1_39P_1_NA_B7));
nor2 N1P_1_179P_1_39P_1_I39_1 (.o(N1P_1_179P_1_39P_1_NA_B3), .i1(N1P_1_179P_1_39P_1_A_B2), .i0(N1P_1_179P_1_39P_1_A_B3));
nor2 N1P_1_179P_1_39P_1_I35_1 (.o(N1P_1_179P_1_39P_1_NA_B1), .i1(N1P_1_179P_1_39P_1_A_B0), .i0(N1P_1_179P_1_39P_1_A_B1));
nor2 N1P_1_179P_1_39P_1_I31_1 (.o(N1P_1_179P_1_39P_1_NA_B7), .i1(N1P_1_179P_1_39P_1_A_B6), .i0(N1P_1_179P_1_39P_1_A_B7));
nor2 N1P_1_179P_1_39P_1_I17_1 (.o(N1P_1_179P_1_39P_1_NA_B5), .i1(N1P_1_179P_1_39P_1_A_B4), .i0(N1P_1_179P_1_39P_1_A_B5));
or5 N1P_1_179P_1_37P_1_I32_1 (.i2(N1P_1_179P_1_37P_1_AB3), .i3(N1P_1_179P_1_37P_1_AB1), .i4(N1P_1_179P_1_37P_1_AG_7), .o(N1P_1_179P_1_UN_1_X74_L85_37P_ALBO), .i1(N1P_1_179P_1_37P_1_AB5), .i0(N1P_1_179P_1_37P_1_AB7));
or5 N1P_1_179P_1_37P_1_I24_1 (.i2(N1P_1_179P_1_37P_1_AB2), .i3(N1P_1_179P_1_37P_1_AB0), .i4(N1P_1_179P_1_37P_1_AL_7), .o(N1P_1_179P_1_UN_1_X74_L85_37P_AGBO), .i1(N1P_1_179P_1_37P_1_AB4), .i0(N1P_1_179P_1_37P_1_AB6));
and2b1 N1P_1_179P_1_37P_1_I41_1 (.o(N1P_1_179P_1_37P_1_A_B0), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I40_1 (.o(N1P_1_179P_1_37P_1_A_B5), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I38_1 (.o(N1P_1_179P_1_37P_1_A_B2), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I37_1 (.o(N1P_1_179P_1_37P_1_A_B7), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I36_1 (.o(N1P_1_179P_1_37P_1_AB6), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I30_1 (.o(N1P_1_179P_1_37P_1_AB7), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I29_1 (.o(N1P_1_179P_1_37P_1_A_B1), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I28_1 (.o(N1P_1_179P_1_37P_1_A_B4), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I26_1 (.o(N1P_1_179P_1_37P_1_A_B6), .i1(XGND), .i0(XGND));
and2b1 N1P_1_179P_1_37P_1_I22_1 (.o(N1P_1_179P_1_37P_1_A_B3), .i1(XGND), .i0(XGND));
and4b1 N1P_1_179P_1_37P_1_I21_1 (.i3(N1P_1_179P_1_37P_1_NA_B5), .i2(XGND), .o(N1P_1_179P_1_37P_1_AB3), .i1(N1P_1_179P_1_37P_1_NA_B7), .i0(XGND));
and4b1 N1P_1_179P_1_37P_1_I20_1 (.i3(N1P_1_179P_1_37P_1_NA_B5), .i2(XGND), .o(N1P_1_179P_1_37P_1_AB2), .i1(N1P_1_179P_1_37P_1_NA_B7), .i0(XGND));
and5b1 N1P_1_179P_1_37P_1_I25_1 (.i4(N1P_1_179P_1_37P_1_NA_B5), .i3(N1P_1_179P_1_37P_1_NA_B3), .i2(XGND), .o(N1P_1_179P_1_37P_1_AB0), .i1(N1P_1_179P_1_37P_1_NA_B7), .i0(XGND));
and5b1 N1P_1_179P_1_37P_1_I16_1 (.i4(N1P_1_179P_1_37P_1_NA_B5), .i3(N1P_1_179P_1_37P_1_NA_B3), .i2(XGND), .o(N1P_1_179P_1_37P_1_AB1), .i1(N1P_1_179P_1_37P_1_NA_B7), .i0(XGND));
and3b1 N1P_1_179P_1_37P_1_I27_1 (.i2(XGND), .o(N1P_1_179P_1_37P_1_AB4), .i1(N1P_1_179P_1_37P_1_NA_B7), .i0(XGND));
and3b1 N1P_1_179P_1_37P_1_I15_1 (.i2(XGND), .o(N1P_1_179P_1_37P_1_AB5), .i1(N1P_1_179P_1_37P_1_NA_B7), .i0(XGND));
and5 N1P_1_179P_1_37P_1_I23_1 (.i2(N1P_1_179P_1_37P_1_NA_B3), .i3(N1P_1_179P_1_37P_1_NA_B1), .i4(XGND), .o(N1P_1_179P_1_37P_1_AEBO), .i1(N1P_1_179P_1_37P_1_NA_B5), .i0(N1P_1_179P_1_37P_1_NA_B7));
and5 N1P_1_179P_1_37P_1_I19_1 (.i2(N1P_1_179P_1_37P_1_NA_B3), .i3(N1P_1_179P_1_37P_1_NA_B1), .i4(N1P_1_LAST_READ[19]), .o(N1P_1_179P_1_37P_1_AL_7), .i1(N1P_1_179P_1_37P_1_NA_B5), .i0(N1P_1_179P_1_37P_1_NA_B7));
and5 N1P_1_179P_1_37P_1_I18_1 (.i2(N1P_1_179P_1_37P_1_NA_B3), .i3(N1P_1_179P_1_37P_1_NA_B1), .i4(N1P_1_LAST_WRITE[19]), .o(N1P_1_179P_1_37P_1_AG_7), .i1(N1P_1_179P_1_37P_1_NA_B5), .i0(N1P_1_179P_1_37P_1_NA_B7));
nor2 N1P_1_179P_1_37P_1_I39_1 (.o(N1P_1_179P_1_37P_1_NA_B3), .i1(N1P_1_179P_1_37P_1_A_B2), .i0(N1P_1_179P_1_37P_1_A_B3));
nor2 N1P_1_179P_1_37P_1_I35_1 (.o(N1P_1_179P_1_37P_1_NA_B1), .i1(N1P_1_179P_1_37P_1_A_B0), .i0(N1P_1_179P_1_37P_1_A_B1));
nor2 N1P_1_179P_1_37P_1_I31_1 (.o(N1P_1_179P_1_37P_1_NA_B7), .i1(N1P_1_179P_1_37P_1_A_B6), .i0(N1P_1_179P_1_37P_1_A_B7));
nor2 N1P_1_179P_1_37P_1_I17_1 (.o(N1P_1_179P_1_37P_1_NA_B5), .i1(N1P_1_179P_1_37P_1_A_B4), .i0(N1P_1_179P_1_37P_1_A_B5));
or5 N1P_1_179P_1_26P_1_I32_1 (.i2(N1P_1_179P_1_26P_1_AB3), .i3(N1P_1_179P_1_26P_1_AB1), .i4(N1P_1_179P_1_26P_1_AG_7), .o(N1P_1_179P_1_UN_1_X74_L85_26P_ALBO), .i1(N1P_1_179P_1_26P_1_AB5), .i0(N1P_1_179P_1_26P_1_AB7));
or5 N1P_1_179P_1_26P_1_I24_1 (.i2(N1P_1_179P_1_26P_1_AB2), .i3(N1P_1_179P_1_26P_1_AB0), .i4(N1P_1_179P_1_26P_1_AL_7), .o(N1P_1_179P_1_UN_1_X74_L85_26P_AGBO), .i1(N1P_1_179P_1_26P_1_AB4), .i0(N1P_1_179P_1_26P_1_AB6));
and2b1 N1P_1_179P_1_26P_1_I41_1 (.o(N1P_1_179P_1_26P_1_A_B0), .i1(N1P_1_LAST_WRITE[15]), .i0(N1P_1_LAST_READ[15]));
and2b1 N1P_1_179P_1_26P_1_I40_1 (.o(N1P_1_179P_1_26P_1_A_B5), .i1(N1P_1_LAST_READ[17]), .i0(N1P_1_LAST_WRITE[17]));
and2b1 N1P_1_179P_1_26P_1_I38_1 (.o(N1P_1_179P_1_26P_1_A_B2), .i1(N1P_1_LAST_WRITE[16]), .i0(N1P_1_LAST_READ[16]));
and2b1 N1P_1_179P_1_26P_1_I37_1 (.o(N1P_1_179P_1_26P_1_A_B7), .i1(N1P_1_LAST_READ[18]), .i0(N1P_1_LAST_WRITE[18]));
and2b1 N1P_1_179P_1_26P_1_I36_1 (.o(N1P_1_179P_1_26P_1_AB6), .i1(N1P_1_LAST_READ[18]), .i0(N1P_1_LAST_WRITE[18]));
and2b1 N1P_1_179P_1_26P_1_I30_1 (.o(N1P_1_179P_1_26P_1_AB7), .i1(N1P_1_LAST_WRITE[18]), .i0(N1P_1_LAST_READ[18]));
and2b1 N1P_1_179P_1_26P_1_I29_1 (.o(N1P_1_179P_1_26P_1_A_B1), .i1(N1P_1_LAST_READ[15]), .i0(N1P_1_LAST_WRITE[15]));
and2b1 N1P_1_179P_1_26P_1_I28_1 (.o(N1P_1_179P_1_26P_1_A_B4), .i1(N1P_1_LAST_WRITE[17]), .i0(N1P_1_LAST_READ[17]));
and2b1 N1P_1_179P_1_26P_1_I26_1 (.o(N1P_1_179P_1_26P_1_A_B6), .i1(N1P_1_LAST_WRITE[18]), .i0(N1P_1_LAST_READ[18]));
and2b1 N1P_1_179P_1_26P_1_I22_1 (.o(N1P_1_179P_1_26P_1_A_B3), .i1(N1P_1_LAST_READ[16]), .i0(N1P_1_LAST_WRITE[16]));
and4b1 N1P_1_179P_1_26P_1_I21_1 (.i3(N1P_1_179P_1_26P_1_NA_B5), .i2(N1P_1_LAST_WRITE[16]), .o(N1P_1_179P_1_26P_1_AB3), .i1(N1P_1_179P_1_26P_1_NA_B7), .i0(N1P_1_LAST_READ[16]));
and4b1 N1P_1_179P_1_26P_1_I20_1 (.i3(N1P_1_179P_1_26P_1_NA_B5), .i2(N1P_1_LAST_READ[16]), .o(N1P_1_179P_1_26P_1_AB2), .i1(N1P_1_179P_1_26P_1_NA_B7), .i0(N1P_1_LAST_WRITE[16]));
and5b1 N1P_1_179P_1_26P_1_I25_1 (.i4(N1P_1_179P_1_26P_1_NA_B5), .i3(N1P_1_179P_1_26P_1_NA_B3), .i2(N1P_1_LAST_READ[15]), .o(N1P_1_179P_1_26P_1_AB0), .i1(N1P_1_179P_1_26P_1_NA_B7), .i0(N1P_1_LAST_WRITE[15]));
and5b1 N1P_1_179P_1_26P_1_I16_1 (.i4(N1P_1_179P_1_26P_1_NA_B5), .i3(N1P_1_179P_1_26P_1_NA_B3), .i2(N1P_1_LAST_WRITE[15]), .o(N1P_1_179P_1_26P_1_AB1), .i1(N1P_1_179P_1_26P_1_NA_B7), .i0(N1P_1_LAST_READ[15]));
and3b1 N1P_1_179P_1_26P_1_I27_1 (.i2(N1P_1_LAST_READ[17]), .o(N1P_1_179P_1_26P_1_AB4), .i1(N1P_1_179P_1_26P_1_NA_B7), .i0(N1P_1_LAST_WRITE[17]));
and3b1 N1P_1_179P_1_26P_1_I15_1 (.i2(N1P_1_LAST_WRITE[17]), .o(N1P_1_179P_1_26P_1_AB5), .i1(N1P_1_179P_1_26P_1_NA_B7), .i0(N1P_1_LAST_READ[17]));
and5 N1P_1_179P_1_26P_1_I23_1 (.i2(N1P_1_179P_1_26P_1_NA_B3), .i3(N1P_1_179P_1_26P_1_NA_B1), .i4(XGND), .o(N1P_1_179P_1_26P_1_AEBO), .i1(N1P_1_179P_1_26P_1_NA_B5), .i0(N1P_1_179P_1_26P_1_NA_B7));
and5 N1P_1_179P_1_26P_1_I19_1 (.i2(N1P_1_179P_1_26P_1_NA_B3), .i3(N1P_1_179P_1_26P_1_NA_B1), .i4(N1P_1_LAST_READ[14]), .o(N1P_1_179P_1_26P_1_AL_7), .i1(N1P_1_179P_1_26P_1_NA_B5), .i0(N1P_1_179P_1_26P_1_NA_B7));
and5 N1P_1_179P_1_26P_1_I18_1 (.i2(N1P_1_179P_1_26P_1_NA_B3), .i3(N1P_1_179P_1_26P_1_NA_B1), .i4(N1P_1_LAST_WRITE[14]), .o(N1P_1_179P_1_26P_1_AG_7), .i1(N1P_1_179P_1_26P_1_NA_B5), .i0(N1P_1_179P_1_26P_1_NA_B7));
nor2 N1P_1_179P_1_26P_1_I39_1 (.o(N1P_1_179P_1_26P_1_NA_B3), .i1(N1P_1_179P_1_26P_1_A_B2), .i0(N1P_1_179P_1_26P_1_A_B3));
nor2 N1P_1_179P_1_26P_1_I35_1 (.o(N1P_1_179P_1_26P_1_NA_B1), .i1(N1P_1_179P_1_26P_1_A_B0), .i0(N1P_1_179P_1_26P_1_A_B1));
nor2 N1P_1_179P_1_26P_1_I31_1 (.o(N1P_1_179P_1_26P_1_NA_B7), .i1(N1P_1_179P_1_26P_1_A_B6), .i0(N1P_1_179P_1_26P_1_A_B7));
nor2 N1P_1_179P_1_26P_1_I17_1 (.o(N1P_1_179P_1_26P_1_NA_B5), .i1(N1P_1_179P_1_26P_1_A_B4), .i0(N1P_1_179P_1_26P_1_A_B5));
or5 N1P_1_179P_1_4P_1_I32_1 (.i2(N1P_1_179P_1_4P_1_AB3), .i3(N1P_1_179P_1_4P_1_AB1), .i4(N1P_1_179P_1_4P_1_AG_7), .o(N1P_1_179P_1_UN_1_X74_L85_39P_B0), .i1(N1P_1_179P_1_4P_1_AB5), .i0(N1P_1_179P_1_4P_1_AB7));
or5 N1P_1_179P_1_4P_1_I24_1 (.i2(N1P_1_179P_1_4P_1_AB2), .i3(N1P_1_179P_1_4P_1_AB0), .i4(N1P_1_179P_1_4P_1_AL_7), .o(N1P_1_179P_1_UN_1_X74_L85_39P_A0), .i1(N1P_1_179P_1_4P_1_AB4), .i0(N1P_1_179P_1_4P_1_AB6));
and2b1 N1P_1_179P_1_4P_1_I41_1 (.o(N1P_1_179P_1_4P_1_A_B0), .i1(N1P_1_LAST_WRITE[5]), .i0(N1P_1_LAST_READ[5]));
and2b1 N1P_1_179P_1_4P_1_I40_1 (.o(N1P_1_179P_1_4P_1_A_B5), .i1(N1P_1_LAST_READ[7]), .i0(N1P_1_LAST_WRITE[7]));
and2b1 N1P_1_179P_1_4P_1_I38_1 (.o(N1P_1_179P_1_4P_1_A_B2), .i1(N1P_1_LAST_WRITE[6]), .i0(N1P_1_LAST_READ[6]));
and2b1 N1P_1_179P_1_4P_1_I37_1 (.o(N1P_1_179P_1_4P_1_A_B7), .i1(N1P_1_LAST_READ[8]), .i0(N1P_1_LAST_WRITE[8]));
and2b1 N1P_1_179P_1_4P_1_I36_1 (.o(N1P_1_179P_1_4P_1_AB6), .i1(N1P_1_LAST_READ[8]), .i0(N1P_1_LAST_WRITE[8]));
and2b1 N1P_1_179P_1_4P_1_I30_1 (.o(N1P_1_179P_1_4P_1_AB7), .i1(N1P_1_LAST_WRITE[8]), .i0(N1P_1_LAST_READ[8]));
and2b1 N1P_1_179P_1_4P_1_I29_1 (.o(N1P_1_179P_1_4P_1_A_B1), .i1(N1P_1_LAST_READ[5]), .i0(N1P_1_LAST_WRITE[5]));
and2b1 N1P_1_179P_1_4P_1_I28_1 (.o(N1P_1_179P_1_4P_1_A_B4), .i1(N1P_1_LAST_WRITE[7]), .i0(N1P_1_LAST_READ[7]));
and2b1 N1P_1_179P_1_4P_1_I26_1 (.o(N1P_1_179P_1_4P_1_A_B6), .i1(N1P_1_LAST_WRITE[8]), .i0(N1P_1_LAST_READ[8]));
and2b1 N1P_1_179P_1_4P_1_I22_1 (.o(N1P_1_179P_1_4P_1_A_B3), .i1(N1P_1_LAST_READ[6]), .i0(N1P_1_LAST_WRITE[6]));
and4b1 N1P_1_179P_1_4P_1_I21_1 (.i3(N1P_1_179P_1_4P_1_NA_B5), .i2(N1P_1_LAST_WRITE[6]), .o(N1P_1_179P_1_4P_1_AB3), .i1(N1P_1_179P_1_4P_1_NA_B7), .i0(N1P_1_LAST_READ[6]));
and4b1 N1P_1_179P_1_4P_1_I20_1 (.i3(N1P_1_179P_1_4P_1_NA_B5), .i2(N1P_1_LAST_READ[6]), .o(N1P_1_179P_1_4P_1_AB2), .i1(N1P_1_179P_1_4P_1_NA_B7), .i0(N1P_1_LAST_WRITE[6]));
and5b1 N1P_1_179P_1_4P_1_I25_1 (.i4(N1P_1_179P_1_4P_1_NA_B5), .i3(N1P_1_179P_1_4P_1_NA_B3), .i2(N1P_1_LAST_READ[5]), .o(N1P_1_179P_1_4P_1_AB0), .i1(N1P_1_179P_1_4P_1_NA_B7), .i0(N1P_1_LAST_WRITE[5]));
and5b1 N1P_1_179P_1_4P_1_I16_1 (.i4(N1P_1_179P_1_4P_1_NA_B5), .i3(N1P_1_179P_1_4P_1_NA_B3), .i2(N1P_1_LAST_WRITE[5]), .o(N1P_1_179P_1_4P_1_AB1), .i1(N1P_1_179P_1_4P_1_NA_B7), .i0(N1P_1_LAST_READ[5]));
and3b1 N1P_1_179P_1_4P_1_I27_1 (.i2(N1P_1_LAST_READ[7]), .o(N1P_1_179P_1_4P_1_AB4), .i1(N1P_1_179P_1_4P_1_NA_B7), .i0(N1P_1_LAST_WRITE[7]));
and3b1 N1P_1_179P_1_4P_1_I15_1 (.i2(N1P_1_LAST_WRITE[7]), .o(N1P_1_179P_1_4P_1_AB5), .i1(N1P_1_179P_1_4P_1_NA_B7), .i0(N1P_1_LAST_READ[7]));
and5 N1P_1_179P_1_4P_1_I23_1 (.i2(N1P_1_179P_1_4P_1_NA_B3), .i3(N1P_1_179P_1_4P_1_NA_B1), .i4(XGND), .o(N1P_1_179P_1_4P_1_AEBO), .i1(N1P_1_179P_1_4P_1_NA_B5), .i0(N1P_1_179P_1_4P_1_NA_B7));
and5 N1P_1_179P_1_4P_1_I19_1 (.i2(N1P_1_179P_1_4P_1_NA_B3), .i3(N1P_1_179P_1_4P_1_NA_B1), .i4(N1P_1_LAST_READ[4]), .o(N1P_1_179P_1_4P_1_AL_7), .i1(N1P_1_179P_1_4P_1_NA_B5), .i0(N1P_1_179P_1_4P_1_NA_B7));
and5 N1P_1_179P_1_4P_1_I18_1 (.i2(N1P_1_179P_1_4P_1_NA_B3), .i3(N1P_1_179P_1_4P_1_NA_B1), .i4(N1P_1_LAST_WRITE[4]), .o(N1P_1_179P_1_4P_1_AG_7), .i1(N1P_1_179P_1_4P_1_NA_B5), .i0(N1P_1_179P_1_4P_1_NA_B7));
nor2 N1P_1_179P_1_4P_1_I39_1 (.o(N1P_1_179P_1_4P_1_NA_B3), .i1(N1P_1_179P_1_4P_1_A_B2), .i0(N1P_1_179P_1_4P_1_A_B3));
nor2 N1P_1_179P_1_4P_1_I35_1 (.o(N1P_1_179P_1_4P_1_NA_B1), .i1(N1P_1_179P_1_4P_1_A_B0), .i0(N1P_1_179P_1_4P_1_A_B1));
nor2 N1P_1_179P_1_4P_1_I31_1 (.o(N1P_1_179P_1_4P_1_NA_B7), .i1(N1P_1_179P_1_4P_1_A_B6), .i0(N1P_1_179P_1_4P_1_A_B7));
nor2 N1P_1_179P_1_4P_1_I17_1 (.o(N1P_1_179P_1_4P_1_NA_B5), .i1(N1P_1_179P_1_4P_1_A_B4), .i0(N1P_1_179P_1_4P_1_A_B5));
or5 N1P_1_179P_1_15P_1_I32_1 (.i2(N1P_1_179P_1_15P_1_AB3), .i3(N1P_1_179P_1_15P_1_AB1), .i4(N1P_1_179P_1_15P_1_AG_7), .o(N1P_1_179P_1_UN_1_X74_L85_15P_ALBO), .i1(N1P_1_179P_1_15P_1_AB5), .i0(N1P_1_179P_1_15P_1_AB7));
or5 N1P_1_179P_1_15P_1_I24_1 (.i2(N1P_1_179P_1_15P_1_AB2), .i3(N1P_1_179P_1_15P_1_AB0), .i4(N1P_1_179P_1_15P_1_AL_7), .o(N1P_1_179P_1_UN_1_X74_L85_15P_AGBO), .i1(N1P_1_179P_1_15P_1_AB4), .i0(N1P_1_179P_1_15P_1_AB6));
and2b1 N1P_1_179P_1_15P_1_I41_1 (.o(N1P_1_179P_1_15P_1_A_B0), .i1(N1P_1_LAST_WRITE[10]), .i0(N1P_1_LAST_READ[10]));
and2b1 N1P_1_179P_1_15P_1_I40_1 (.o(N1P_1_179P_1_15P_1_A_B5), .i1(N1P_1_LAST_READ[12]), .i0(N1P_1_LAST_WRITE[12]));
and2b1 N1P_1_179P_1_15P_1_I38_1 (.o(N1P_1_179P_1_15P_1_A_B2), .i1(N1P_1_LAST_WRITE[11]), .i0(N1P_1_LAST_READ[11]));
and2b1 N1P_1_179P_1_15P_1_I37_1 (.o(N1P_1_179P_1_15P_1_A_B7), .i1(N1P_1_LAST_READ[13]), .i0(N1P_1_LAST_WRITE[13]));
and2b1 N1P_1_179P_1_15P_1_I36_1 (.o(N1P_1_179P_1_15P_1_AB6), .i1(N1P_1_LAST_READ[13]), .i0(N1P_1_LAST_WRITE[13]));
and2b1 N1P_1_179P_1_15P_1_I30_1 (.o(N1P_1_179P_1_15P_1_AB7), .i1(N1P_1_LAST_WRITE[13]), .i0(N1P_1_LAST_READ[13]));
and2b1 N1P_1_179P_1_15P_1_I29_1 (.o(N1P_1_179P_1_15P_1_A_B1), .i1(N1P_1_LAST_READ[10]), .i0(N1P_1_LAST_WRITE[10]));
and2b1 N1P_1_179P_1_15P_1_I28_1 (.o(N1P_1_179P_1_15P_1_A_B4), .i1(N1P_1_LAST_WRITE[12]), .i0(N1P_1_LAST_READ[12]));
and2b1 N1P_1_179P_1_15P_1_I26_1 (.o(N1P_1_179P_1_15P_1_A_B6), .i1(N1P_1_LAST_WRITE[13]), .i0(N1P_1_LAST_READ[13]));
and2b1 N1P_1_179P_1_15P_1_I22_1 (.o(N1P_1_179P_1_15P_1_A_B3), .i1(N1P_1_LAST_READ[11]), .i0(N1P_1_LAST_WRITE[11]));
and4b1 N1P_1_179P_1_15P_1_I21_1 (.i3(N1P_1_179P_1_15P_1_NA_B5), .i2(N1P_1_LAST_WRITE[11]), .o(N1P_1_179P_1_15P_1_AB3), .i1(N1P_1_179P_1_15P_1_NA_B7), .i0(N1P_1_LAST_READ[11]));
and4b1 N1P_1_179P_1_15P_1_I20_1 (.i3(N1P_1_179P_1_15P_1_NA_B5), .i2(N1P_1_LAST_READ[11]), .o(N1P_1_179P_1_15P_1_AB2), .i1(N1P_1_179P_1_15P_1_NA_B7), .i0(N1P_1_LAST_WRITE[11]));
and5b1 N1P_1_179P_1_15P_1_I25_1 (.i4(N1P_1_179P_1_15P_1_NA_B5), .i3(N1P_1_179P_1_15P_1_NA_B3), .i2(N1P_1_LAST_READ[10]), .o(N1P_1_179P_1_15P_1_AB0), .i1(N1P_1_179P_1_15P_1_NA_B7), .i0(N1P_1_LAST_WRITE[10]));
and5b1 N1P_1_179P_1_15P_1_I16_1 (.i4(N1P_1_179P_1_15P_1_NA_B5), .i3(N1P_1_179P_1_15P_1_NA_B3), .i2(N1P_1_LAST_WRITE[10]), .o(N1P_1_179P_1_15P_1_AB1), .i1(N1P_1_179P_1_15P_1_NA_B7), .i0(N1P_1_LAST_READ[10]));
and3b1 N1P_1_179P_1_15P_1_I27_1 (.i2(N1P_1_LAST_READ[12]), .o(N1P_1_179P_1_15P_1_AB4), .i1(N1P_1_179P_1_15P_1_NA_B7), .i0(N1P_1_LAST_WRITE[12]));
and3b1 N1P_1_179P_1_15P_1_I15_1 (.i2(N1P_1_LAST_WRITE[12]), .o(N1P_1_179P_1_15P_1_AB5), .i1(N1P_1_179P_1_15P_1_NA_B7), .i0(N1P_1_LAST_READ[12]));
and5 N1P_1_179P_1_15P_1_I23_1 (.i2(N1P_1_179P_1_15P_1_NA_B3), .i3(N1P_1_179P_1_15P_1_NA_B1), .i4(XGND), .o(N1P_1_179P_1_15P_1_AEBO), .i1(N1P_1_179P_1_15P_1_NA_B5), .i0(N1P_1_179P_1_15P_1_NA_B7));
and5 N1P_1_179P_1_15P_1_I19_1 (.i2(N1P_1_179P_1_15P_1_NA_B3), .i3(N1P_1_179P_1_15P_1_NA_B1), .i4(N1P_1_LAST_READ[9]), .o(N1P_1_179P_1_15P_1_AL_7), .i1(N1P_1_179P_1_15P_1_NA_B5), .i0(N1P_1_179P_1_15P_1_NA_B7));
and5 N1P_1_179P_1_15P_1_I18_1 (.i2(N1P_1_179P_1_15P_1_NA_B3), .i3(N1P_1_179P_1_15P_1_NA_B1), .i4(N1P_1_LAST_WRITE[9]), .o(N1P_1_179P_1_15P_1_AG_7), .i1(N1P_1_179P_1_15P_1_NA_B5), .i0(N1P_1_179P_1_15P_1_NA_B7));
nor2 N1P_1_179P_1_15P_1_I39_1 (.o(N1P_1_179P_1_15P_1_NA_B3), .i1(N1P_1_179P_1_15P_1_A_B2), .i0(N1P_1_179P_1_15P_1_A_B3));
nor2 N1P_1_179P_1_15P_1_I35_1 (.o(N1P_1_179P_1_15P_1_NA_B1), .i1(N1P_1_179P_1_15P_1_A_B0), .i0(N1P_1_179P_1_15P_1_A_B1));
nor2 N1P_1_179P_1_15P_1_I31_1 (.o(N1P_1_179P_1_15P_1_NA_B7), .i1(N1P_1_179P_1_15P_1_A_B6), .i0(N1P_1_179P_1_15P_1_A_B7));
nor2 N1P_1_179P_1_15P_1_I17_1 (.o(N1P_1_179P_1_15P_1_NA_B5), .i1(N1P_1_179P_1_15P_1_A_B4), .i0(N1P_1_179P_1_15P_1_A_B5));
and5 N1P_1_179P_1_2P_1 (.i2(N1P_1_179P_1_UN_1_AND5_2P_I2), .i3(N1P_1_179P_1_UN_1_AND5_2P_I3), .i4(N1P_1_179P_1_UN_1_AND5_2P_I4), .o(N1P_1_179P_1_UN_1_AND2_41P_I1), .i1(N1P_1_179P_1_UN_1_AND5_2P_I1), .i0(N1P_1_179P_1_UN_1_AND5_2P_I0));
and2 N1P_1_179P_1_42P_1 (.o(BREAD_EN_n), .i1(N1P_1_179P_1_UN_1_AND2_41P_I1), .i0(N1P_1_179P_1_UN_1_AND2_42P_I0));
and2 N1P_1_179P_1_41P_1 (.o(BWRITE_EN_n), .i1(N1P_1_179P_1_UN_1_AND2_41P_I1), .i0(N1P_1_179P_1_UN_1_AND2_41P_I0));
or2 N1P_1_179P_1_40P_1 (.o(N1P_1_179P_1_UN_1_AND2_42P_I0), .i1(N1P_1_179P_1_UN_1_OR2_40P_I1), .i0(N1P_1_179P_1_UN_1_OR2_40P_I0));
inv N1P_1_181P_1 (.i(FIFO_RESET_n), .o(N1P_1_FIFO_RESET));
inv N1P_1_172P_1 (.i(SEL2_n), .o(N1P_1_SEL2));
inv N1P_1_170P_1 (.i(SEL1_n), .o(N1P_1_SEL1));
nand2 N75P_1 (.o(MEMACK2_n), .i1(MDTACK), .i0(SEL2));
nand2 N58P_1 (.o(MEMACK1_n), .i1(MDTACK), .i0(SEL1));
and2 N54P_1 (.o(REQ1_n), .i1(UN_1_AND2_54P_I1), .i0(UN_1_AND2_54P_I0));
nor2 N51P_1 (.o(UN_1_NOR2_50P_I0), .i1(MDTACK), .i0(BRW_n));
nor2 N50P_1 (.o(MEM_WRITE_ENABLE_n), .i1(SEL2), .i0(UN_1_NOR2_50P_I0));
or2 N67P_1 (.o(READ_BLKACK_n), .i1(UN_1_INV_66P_O), .i0(MEMACK1_n));
or2 N55P_1 (.o(UN_1_AND2_54P_I1), .i1(BREAD_EN_n), .i0(MEMREQ1_n));
or2 N53P_1 (.o(REQ2_IN_n), .i1(BWRITE_EN_n), .i0(MEMREQ2_n));
or2 N46P_1 (.o(UN_1_AND2_54P_I0), .i1(MEMREQ1_n), .i0(TESTMEM2_n));
or2 N45P_1 (.o(MEMREQ1_n), .i1(MODSEL_n), .i0(MEMSPACE_n));
inv N76P_1 (.i(SIMM_EN_[0]), .o(UN_1_FDC_65P_CLR));
inv N74P_1 (.i(SIMM_EN_[5]), .o(UN_1_FDC_65P_C));
inv N68P_1 (.i(MEMREQ1_n), .o(MEMREQ1));
inv N66P_1 (.i(UN_1_FDC_65P_Q), .o(UN_1_INV_66P_O));
inv N60P_1 (.i(SEL1_n), .o(SEL1));
inv N59P_1 (.i(REQ1_n), .o(REQ1));
inv N52P_1 (.i(SEL2_n), .o(SEL2));
inv N44P_1 (.i(TESTMEM2), .o(TESTMEM2_n));
obuf N2P_1_8 (.i(SIMM_EN_[7]), .o(XSIMM_EN_[7]));
obuf N2P_1_7 (.o(XSIMM_EN_[6]), .i(SIMM_EN_[6]));
obuf N2P_1_6 (.o(XSIMM_EN_[5]), .i(SIMM_EN_[5]));
obuf N2P_1_5 (.o(XSIMM_EN_[4]), .i(SIMM_EN_[4]));
obuf N2P_1_4 (.o(XSIMM_EN_[3]), .i(SIMM_EN_[3]));
obuf N2P_1_3 (.o(XSIMM_EN_[2]), .i(SIMM_EN_[2]));
obuf N2P_1_2 (.o(XSIMM_EN_[1]), .i(SIMM_EN_[1]));
obuf N2P_1_1 (.o(XSIMM_EN_[0]), .i(SIMM_EN_[0]));
obuf N84P_1_5 (.i(UN_1_IBUF_82P_O[4]), .o(SPARES[4]));
obuf N84P_1_4 (.o(SPARES[3]), .i(UN_1_IBUF_82P_O[3]));
obuf N84P_1_3 (.o(SPARES[2]), .i(UN_1_IBUF_82P_O[2]));
obuf N84P_1_2 (.o(SPARES[1]), .i(UN_1_IBUF_82P_O[1]));
obuf N84P_1_1 (.o(SPARES[0]), .i(UN_1_IBUF_82P_O[0]));
obuf N7P_1_20 (.i(BWR_ADD[21]), .o(XBWR_ADD[21]));
obuf N7P_1_19 (.o(XBWR_ADD[20]), .i(BWR_ADD[20]));
obuf N7P_1_18 (.o(XBWR_ADD[19]), .i(BWR_ADD[19]));
obuf N7P_1_17 (.o(XBWR_ADD[18]), .i(BWR_ADD[18]));
obuf N7P_1_16 (.o(XBWR_ADD[17]), .i(BWR_ADD[17]));
obuf N7P_1_15 (.o(XBWR_ADD[16]), .i(BWR_ADD[16]));
obuf N7P_1_14 (.o(XBWR_ADD[15]), .i(BWR_ADD[15]));
obuf N7P_1_13 (.o(XBWR_ADD[14]), .i(BWR_ADD[14]));
obuf N7P_1_12 (.o(XBWR_ADD[13]), .i(BWR_ADD[13]));
obuf N7P_1_11 (.o(XBWR_ADD[12]), .i(BWR_ADD[12]));
obuf N7P_1_10 (.o(XBWR_ADD[11]), .i(BWR_ADD[11]));
obuf N7P_1_9 (.o(XBWR_ADD[10]), .i(BWR_ADD[10]));
obuf N7P_1_8 (.o(XBWR_ADD[9]), .i(BWR_ADD[9]));
obuf N7P_1_7 (.o(XBWR_ADD[8]), .i(BWR_ADD[8]));
obuf N7P_1_6 (.o(XBWR_ADD[7]), .i(BWR_ADD[7]));
obuf N7P_1_5 (.o(XBWR_ADD[6]), .i(BWR_ADD[6]));
obuf N7P_1_4 (.o(XBWR_ADD[5]), .i(BWR_ADD[5]));
obuf N7P_1_3 (.o(XBWR_ADD[4]), .i(BWR_ADD[4]));
obuf N7P_1_2 (.o(XBWR_ADD[3]), .i(BWR_ADD[3]));
obuf N7P_1_1 (.o(XBWR_ADD[2]), .i(BWR_ADD[2]));
obuf N85P_1 (.i(UN_1_IBUF_83P_O), .o(SDOUT));
obuf N79P_1 (.i(XVDD), .o(M2));
obuf N3P_1 (.i(MEM_WRITE_ENABLE_n), .o(XMEM_WRITE_ENABLE_n));
obuf N4P_1 (.i(MEMACK1_n), .o(XMEMACK1_n));
obuf N5P_1 (.i(MEMACK2_n), .o(XMEMACK2_n));
obuf N8P_1 (.i(REQ2_n), .o(XREQ2_n));
obuf N9P_1 (.i(REQ1_n), .o(XREQ1_n));
ibuf N82P_1_5 (.i(SPARES[9]), .o(UN_1_IBUF_82P_O[4]));
ibuf N82P_1_4 (.o(UN_1_IBUF_82P_O[3]), .i(SPARES[8]));
ibuf N82P_1_3 (.o(UN_1_IBUF_82P_O[2]), .i(SPARES[7]));
ibuf N82P_1_2 (.o(UN_1_IBUF_82P_O[1]), .i(SPARES[6]));
ibuf N82P_1_1 (.o(UN_1_IBUF_82P_O[0]), .i(SPARES[5]));
ibuf N29P_1_23 (.i(XBBA[24]), .o(BBA[24]));
ibuf N29P_1_22 (.o(BBA[23]), .i(XBBA[23]));
ibuf N29P_1_21 (.o(BBA[22]), .i(XBBA[22]));
ibuf N29P_1_20 (.o(BBA[21]), .i(XBBA[21]));
ibuf N29P_1_19 (.o(BBA[20]), .i(XBBA[20]));
ibuf N29P_1_18 (.o(BBA[19]), .i(XBBA[19]));
ibuf N29P_1_17 (.o(BBA[18]), .i(XBBA[18]));
ibuf N29P_1_16 (.o(BBA[17]), .i(XBBA[17]));
ibuf N29P_1_15 (.o(BBA[16]), .i(XBBA[16]));
ibuf N29P_1_14 (.o(BBA[15]), .i(XBBA[15]));
ibuf N29P_1_13 (.o(BBA[14]), .i(XBBA[14]));
ibuf N29P_1_12 (.o(BBA[13]), .i(XBBA[13]));
ibuf N29P_1_11 (.o(BBA[12]), .i(XBBA[12]));
ibuf N29P_1_10 (.o(BBA[11]), .i(XBBA[11]));
ibuf N29P_1_9 (.o(BBA[10]), .i(XBBA[10]));
ibuf N29P_1_8 (.o(BBA[9]), .i(XBBA[9]));
ibuf N29P_1_7 (.o(BBA[8]), .i(XBBA[8]));
ibuf N29P_1_6 (.o(BBA[7]), .i(XBBA[7]));
ibuf N29P_1_5 (.o(BBA[6]), .i(XBBA[6]));
ibuf N29P_1_4 (.o(BBA[5]), .i(XBBA[5]));
ibuf N29P_1_3 (.o(BBA[4]), .i(XBBA[4]));
ibuf N29P_1_2 (.o(BBA[3]), .i(XBBA[3]));
ibuf N29P_1_1 (.o(BBA[2]), .i(XBBA[2]));
ibuf N83P_1 (.i(SDIN), .o(UN_1_IBUF_83P_O));
ibuf N28P_1 (.i(XSEL1_n), .o(SEL1_n));
ibuf N27P_1 (.i(XSEL2_n), .o(SEL2_n));
ibuf N26P_1 (.i(XFIFO_RESET_n), .o(FIFO_RESET_n));
ibuf N25P_1 (.i(XTESTMEM1), .o(TESTMEM1));
ibuf N24P_1 (.i(XMODSEL_n), .o(MODSEL_n));
ibuf N23P_1 (.i(XMEMSPACE_n), .o(MEMSPACE_n));
ibuf N22P_1 (.i(XTESTMEM2), .o(TESTMEM2));
ibuf N21P_1 (.i(XMEMREQ2_n), .o(MEMREQ2_n));
ibuf N20P_1 (.i(XBRW_n), .o(BRW_n));
ibuf N18P_1 (.i(XMDTACK), .o(MDTACK));
endmodule
`uselib

module xmemfifo_globals();

wire GR;
endmodule

