/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from bregs96t.xcd on Sat Jun  1 12:40:55 1996 */
/* PART 3020PC84-70 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module bregs96t
(SPAREOUT, SPAREIN, M2, DOUT, DIN, BTESTMODE1, BSQCREG_REQ, BSBSELECT, BSBREAD_n, BREG32_63_WR_n, BREG32_63_RD_n, BREGSPACE, BREG_WR_, BREG_RD_, BFIFOREG_WR_n, BFIFOREG_RD_n, BDTACK_REQ_n, BCREG_REG_n, BA, PWRDWN_n, RDATA_n, RTRIG, RESET_n, PROGRAM_n, CCLK);
   output [1:0] SPAREOUT;
   input [1:0] SPAREIN;
   output M2;
   output DOUT;
   input DIN;
   input BTESTMODE1;
   output BSQCREG_REQ;
   input BSBSELECT;
   input BSBREAD_n;
   output BREG32_63_WR_n;
   output BREG32_63_RD_n;
   input BREGSPACE;
   output [15:0] BREG_WR_;
   output [15:0] BREG_RD_;
   output BFIFOREG_WR_n;
   output BFIFOREG_RD_n;
   output BDTACK_REQ_n;
   output BCREG_REG_n;
   input [10:2] BA;
   input PWRDWN_n;
   output RDATA_n;
   input RTRIG;
   input RESET_n;
   input PROGRAM_n;
   input CCLK;
wire [0:0] N92P_2_I35;
wire [1:0] UN_3_AND2_3P_O;
wire [1:0] UN_3_AND2_3P_I0;
wire [15:0] REG_WR_;
wire [15:0] REG_RD_;
wire [10:2] A;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/preprod_board/fec32m/develop/bregs96t/verilog_lib/bregs96t.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

and4 N92P_2_I11_1 (.o(UN_2_AND6_92P_O), .i1(UN_2_AND6_92P_I1), .i0(UN_2_AND6_92P_I0), .i2(UN_2_AND6_92P_I2), .i3(N92P_2_I35[0]));
and3 N92P_2_I8_1 (.o(N92P_2_I35[0]), .i1(UN_2_AND6_92P_I4), .i0(UN_2_AND6_92P_I3), .i2(D_REGSEL));
nand5b4 N265P_1_I40_1 (.o(REG_RD_[0]), .i3(A[4]), .i2(A[5]), .i1(A[3]), .i0(A[2]), .i4(N265P_1_UN_1_NAND5_I34_I4));
nand5 N265P_1_I34_1 (.o(REG_RD_[15]), .i1(A[4]), .i0(A[5]), .i2(A[3]), .i3(A[2]), .i4(N265P_1_UN_1_NAND5_I34_I4));
nand5b2 N265P_1_I39_1 (.o(REG_RD_[10]), .i1(A[4]), .i0(A[2]), .i4(N265P_1_UN_1_NAND5_I34_I4), .i3(A[5]), .i2(A[3]));
nand5b2 N265P_1_I37_1 (.o(REG_RD_[6]), .i1(A[2]), .i0(A[5]), .i4(N265P_1_UN_1_NAND5_I34_I4), .i3(A[4]), .i2(A[3]));
nand5b2 N265P_1_I36_1 (.o(REG_RD_[5]), .i1(A[3]), .i0(A[5]), .i4(N265P_1_UN_1_NAND5_I34_I4), .i3(A[4]), .i2(A[2]));
nand5b2 N265P_1_I32_1 (.o(REG_RD_[9]), .i1(A[4]), .i0(A[3]), .i4(N265P_1_UN_1_NAND5_I34_I4), .i3(A[5]), .i2(A[2]));
nand5b2 N265P_1_I31_1 (.o(REG_RD_[12]), .i1(A[3]), .i0(A[2]), .i4(N265P_1_UN_1_NAND5_I34_I4), .i3(A[5]), .i2(A[4]));
nand5b2 N265P_1_I30_1 (.o(REG_RD_[3]), .i1(A[5]), .i0(A[4]), .i4(N265P_1_UN_1_NAND5_I34_I4), .i3(A[2]), .i2(A[3]));
nand5b3 N265P_1_I38_1 (.o(REG_RD_[4]), .i2(A[3]), .i1(A[2]), .i0(A[5]), .i4(A[4]), .i3(N265P_1_UN_1_NAND5_I34_I4));
nand5b3 N265P_1_I35_1 (.o(REG_RD_[8]), .i2(A[3]), .i1(A[2]), .i0(A[4]), .i4(A[5]), .i3(N265P_1_UN_1_NAND5_I34_I4));
nand5b3 N265P_1_I27_1 (.o(REG_RD_[1]), .i2(A[4]), .i1(A[3]), .i0(A[5]), .i4(A[2]), .i3(N265P_1_UN_1_NAND5_I34_I4));
nand5b3 N265P_1_I26_1 (.o(REG_RD_[2]), .i2(A[5]), .i1(A[2]), .i0(A[4]), .i4(A[3]), .i3(N265P_1_UN_1_NAND5_I34_I4));
nand5b1 N265P_1_I41_1 (.o(REG_RD_[7]), .i4(A[4]), .i0(A[5]), .i3(A[3]), .i2(A[2]), .i1(N265P_1_UN_1_NAND5_I34_I4));
nand5b1 N265P_1_I33_1 (.o(REG_RD_[11]), .i4(A[2]), .i0(A[4]), .i3(A[3]), .i2(A[5]), .i1(N265P_1_UN_1_NAND5_I34_I4));
nand5b1 N265P_1_I29_1 (.o(REG_RD_[13]), .i4(A[2]), .i0(A[3]), .i3(A[4]), .i2(A[5]), .i1(N265P_1_UN_1_NAND5_I34_I4));
nand5b1 N265P_1_I25_1 (.o(REG_RD_[14]), .i4(A[3]), .i0(A[2]), .i3(A[4]), .i2(A[5]), .i1(N265P_1_UN_1_NAND5_I34_I4));
nor2 N265P_1_I28_1 (.o(N265P_1_UN_1_NAND5_I34_I4), .i1(D_REGSEL_n), .i0(REG0_31RD_n));
nand5b4 N264P_1_I40_1 (.o(REG_WR_[0]), .i3(UN_1_4_MERGE_340P_B), .i2(UN_1_4_MERGE_340P_A), .i1(UN_1_4_MERGE_340P_C), .i0(UN_1_4_MERGE_340P_D), .i4(N264P_1_UN_1_NAND5_I34_I4));
nand5 N264P_1_I34_1 (.o(REG_WR_[15]), .i1(UN_1_4_MERGE_340P_B), .i0(UN_1_4_MERGE_340P_A), .i2(UN_1_4_MERGE_340P_C), .i3(UN_1_4_MERGE_340P_D), .i4(N264P_1_UN_1_NAND5_I34_I4));
nand5b2 N264P_1_I39_1 (.o(REG_WR_[10]), .i1(UN_1_4_MERGE_340P_B), .i0(UN_1_4_MERGE_340P_D), .i4(N264P_1_UN_1_NAND5_I34_I4), .i3(UN_1_4_MERGE_340P_A), .i2(UN_1_4_MERGE_340P_C));
nand5b2 N264P_1_I37_1 (.o(REG_WR_[6]), .i1(UN_1_4_MERGE_340P_D), .i0(UN_1_4_MERGE_340P_A), .i4(N264P_1_UN_1_NAND5_I34_I4), .i3(UN_1_4_MERGE_340P_B), .i2(UN_1_4_MERGE_340P_C));
nand5b2 N264P_1_I36_1 (.o(REG_WR_[5]), .i1(UN_1_4_MERGE_340P_C), .i0(UN_1_4_MERGE_340P_A), .i4(N264P_1_UN_1_NAND5_I34_I4), .i3(UN_1_4_MERGE_340P_B), .i2(UN_1_4_MERGE_340P_D));
nand5b2 N264P_1_I32_1 (.o(REG_WR_[9]), .i1(UN_1_4_MERGE_340P_B), .i0(UN_1_4_MERGE_340P_C), .i4(N264P_1_UN_1_NAND5_I34_I4), .i3(UN_1_4_MERGE_340P_A), .i2(UN_1_4_MERGE_340P_D));
nand5b2 N264P_1_I31_1 (.o(REG_WR_[12]), .i1(UN_1_4_MERGE_340P_C), .i0(UN_1_4_MERGE_340P_D), .i4(N264P_1_UN_1_NAND5_I34_I4), .i3(UN_1_4_MERGE_340P_A), .i2(UN_1_4_MERGE_340P_B));
nand5b2 N264P_1_I30_1 (.o(REG_WR_[3]), .i1(UN_1_4_MERGE_340P_A), .i0(UN_1_4_MERGE_340P_B), .i4(N264P_1_UN_1_NAND5_I34_I4), .i3(UN_1_4_MERGE_340P_D), .i2(UN_1_4_MERGE_340P_C));
nand5b3 N264P_1_I38_1 (.o(UN_1_INV_348P_I), .i2(UN_1_4_MERGE_340P_C), .i1(UN_1_4_MERGE_340P_D), .i0(UN_1_4_MERGE_340P_A), .i4(UN_1_4_MERGE_340P_B), .i3(N264P_1_UN_1_NAND5_I34_I4));
nand5b3 N264P_1_I35_1 (.o(REG_WR_[8]), .i2(UN_1_4_MERGE_340P_C), .i1(UN_1_4_MERGE_340P_D), .i0(UN_1_4_MERGE_340P_B), .i4(UN_1_4_MERGE_340P_A), .i3(N264P_1_UN_1_NAND5_I34_I4));
nand5b3 N264P_1_I27_1 (.o(REG_WR_[1]), .i2(UN_1_4_MERGE_340P_B), .i1(UN_1_4_MERGE_340P_C), .i0(UN_1_4_MERGE_340P_A), .i4(UN_1_4_MERGE_340P_D), .i3(N264P_1_UN_1_NAND5_I34_I4));
nand5b3 N264P_1_I26_1 (.o(REG_WR_[2]), .i2(UN_1_4_MERGE_340P_A), .i1(UN_1_4_MERGE_340P_D), .i0(UN_1_4_MERGE_340P_B), .i4(UN_1_4_MERGE_340P_C), .i3(N264P_1_UN_1_NAND5_I34_I4));
nand5b1 N264P_1_I41_1 (.o(REG_WR_[7]), .i4(UN_1_4_MERGE_340P_B), .i0(UN_1_4_MERGE_340P_A), .i3(UN_1_4_MERGE_340P_C), .i2(UN_1_4_MERGE_340P_D), .i1(N264P_1_UN_1_NAND5_I34_I4));
nand5b1 N264P_1_I33_1 (.o(UN_1_INV_346P_I), .i4(UN_1_4_MERGE_340P_D), .i0(UN_1_4_MERGE_340P_B), .i3(UN_1_4_MERGE_340P_C), .i2(UN_1_4_MERGE_340P_A), .i1(N264P_1_UN_1_NAND5_I34_I4));
nand5b1 N264P_1_I29_1 (.o(REG_WR_[13]), .i4(UN_1_4_MERGE_340P_D), .i0(UN_1_4_MERGE_340P_C), .i3(UN_1_4_MERGE_340P_B), .i2(UN_1_4_MERGE_340P_A), .i1(N264P_1_UN_1_NAND5_I34_I4));
nand5b1 N264P_1_I25_1 (.o(REG_WR_[14]), .i4(UN_1_4_MERGE_340P_C), .i0(UN_1_4_MERGE_340P_D), .i3(UN_1_4_MERGE_340P_B), .i2(UN_1_4_MERGE_340P_A), .i1(N264P_1_UN_1_NAND5_I34_I4));
nor2 N264P_1_I28_1 (.o(N264P_1_UN_1_NAND5_I34_I4), .i1(D_REGSEL_n), .i0(REG0_15WR_n));
and2b1 N338P_1 (.o(SQCREG_REQ), .i1(UN_1_AND2_53P_O), .i0(TESTMODE1));
buff N342P_1_4 (.o(UN_1_4_MERGE_340P_A), .i(A[5]));
buff N342P_1_3 (.i(A[4]), .o(UN_1_4_MERGE_340P_B));
buff N342P_1_2 (.i(A[3]), .o(UN_1_4_MERGE_340P_C));
buff N342P_1_1 (.i(A[2]), .o(UN_1_4_MERGE_340P_D));
ibuf N299P_1_9 (.o(A[10]), .i(BA[10]));
ibuf N299P_1_8 (.i(BA[9]), .o(A[9]));
ibuf N299P_1_7 (.i(BA[8]), .o(A[8]));
ibuf N299P_1_6 (.i(BA[7]), .o(A[7]));
ibuf N299P_1_5 (.i(BA[6]), .o(A[6]));
ibuf N299P_1_4 (.i(BA[5]), .o(A[5]));
ibuf N299P_1_3 (.i(BA[4]), .o(A[4]));
ibuf N299P_1_2 (.i(BA[3]), .o(A[3]));
ibuf N299P_1_1 (.i(BA[2]), .o(A[2]));
ibuf N325P_1 (.o(SBSELECT), .i(BSBSELECT));
ibuf N324P_1 (.o(REGSPACE), .i(BREGSPACE));
ibuf N323P_1 (.o(SBREAD_n), .i(BSBREAD_n));
ibuf N293P_1 (.o(TESTMODE1), .i(BTESTMODE1));
ibuf N4P_3_2 (.o(UN_3_AND2_3P_I0[1]), .i(SPAREIN[1]));
ibuf N4P_3_1 (.i(SPAREIN[0]), .o(UN_3_AND2_3P_I0[0]));
ibuf N7P_3 (.o(UN_3_AND2_10P_I0), .i(DIN));
obuf N71P_2 (.o(BDTACK_REQ_n), .i(DTACK_REQ_n));
obuf N285P_1 (.o(BCREG_REG_n), .i(CREG_REG_n));
obuf N296P_1_16 (.o(BREG_RD_[15]), .i(REG_RD_[15]));
obuf N296P_1_15 (.i(REG_RD_[14]), .o(BREG_RD_[14]));
obuf N296P_1_14 (.i(REG_RD_[13]), .o(BREG_RD_[13]));
obuf N296P_1_13 (.i(REG_RD_[12]), .o(BREG_RD_[12]));
obuf N296P_1_12 (.i(REG_RD_[11]), .o(BREG_RD_[11]));
obuf N296P_1_11 (.i(REG_RD_[10]), .o(BREG_RD_[10]));
obuf N296P_1_10 (.i(REG_RD_[9]), .o(BREG_RD_[9]));
obuf N296P_1_9 (.i(REG_RD_[8]), .o(BREG_RD_[8]));
obuf N296P_1_8 (.i(REG_RD_[7]), .o(BREG_RD_[7]));
obuf N296P_1_7 (.i(REG_RD_[6]), .o(BREG_RD_[6]));
obuf N296P_1_6 (.i(REG_RD_[5]), .o(BREG_RD_[5]));
obuf N296P_1_5 (.i(REG_RD_[4]), .o(BREG_RD_[4]));
obuf N296P_1_4 (.i(REG_RD_[3]), .o(BREG_RD_[3]));
obuf N296P_1_3 (.i(REG_RD_[2]), .o(BREG_RD_[2]));
obuf N296P_1_2 (.i(REG_RD_[1]), .o(BREG_RD_[1]));
obuf N296P_1_1 (.i(REG_RD_[0]), .o(BREG_RD_[0]));
obuf N295P_1_16 (.o(BREG_WR_[15]), .i(REG_WR_[15]));
obuf N295P_1_15 (.i(REG_WR_[14]), .o(BREG_WR_[14]));
obuf N295P_1_14 (.i(REG_WR_[13]), .o(BREG_WR_[13]));
obuf N295P_1_13 (.i(REG_WR_[12]), .o(BREG_WR_[12]));
obuf N295P_1_12 (.i(REG_WR_[11]), .o(BREG_WR_[11]));
obuf N295P_1_11 (.i(REG_WR_[10]), .o(BREG_WR_[10]));
obuf N295P_1_10 (.i(REG_WR_[9]), .o(BREG_WR_[9]));
obuf N295P_1_9 (.i(REG_WR_[8]), .o(BREG_WR_[8]));
obuf N295P_1_8 (.i(REG_WR_[7]), .o(BREG_WR_[7]));
obuf N295P_1_7 (.i(REG_WR_[6]), .o(BREG_WR_[6]));
obuf N295P_1_6 (.i(REG_WR_[5]), .o(BREG_WR_[5]));
obuf N295P_1_5 (.i(REG_WR_[4]), .o(BREG_WR_[4]));
obuf N295P_1_4 (.i(REG_WR_[3]), .o(BREG_WR_[3]));
obuf N295P_1_3 (.i(REG_WR_[2]), .o(BREG_WR_[2]));
obuf N295P_1_2 (.i(REG_WR_[1]), .o(BREG_WR_[1]));
obuf N295P_1_1 (.i(REG_WR_[0]), .o(BREG_WR_[0]));
obuf N1P_3_2 (.o(SPAREOUT[1]), .i(UN_3_AND2_3P_O[1]));
obuf N1P_3_1 (.i(UN_3_AND2_3P_O[0]), .o(SPAREOUT[0]));
obuf N11P_3 (.o(M2), .i(XVDD));
obuf N9P_3 (.o(DOUT), .i(UN_3_AND2_10P_O));
obuf N87P_2 (.o(BFIFOREG_WR_n), .i(FIFOREG_WR_n));
obuf N86P_2 (.o(BFIFOREG_RD_n), .i(FIFOREG_RD_n));
obuf N337P_1 (.o(BSQCREG_REQ), .i(SQCREG_REQ));
obuf N334P_1 (.o(BREG32_63_WR_n), .i(REG32_63_WR_n));
obuf N333P_1 (.o(BREG32_63_RD_n), .i(REG32_63_RD_n));
nor2 N283P_1 (.o(UN_1_AND2_232P_I1), .i1(UN_1_NOR2_283P_I1), .i0(UN_1_NOR2_283P_I0));
nand3 N243P_1 (.o(REG32_63_WR_n), .i1(UN_1_INV_234P_O), .i0(REG32_63), .i2(SBREAD_n));
nand3 N242P_1 (.o(REG32_63_RD_n), .i1(UN_1_INV_234P_O), .i0(REG32_63), .i2(SBREAD));
and2 N10P_3 (.o(UN_3_AND2_10P_O), .i1(UN_3_AND2_10P_I0), .i0(UN_3_AND2_10P_I0));
and2 N60P_2 (.o(FIFOREG_REQ), .i1(FIFO_REG), .i0(REG32_63));
and2 N63P_1 (.o(REGSEL), .i1(SBSELECT), .i0(REGSPACE));
and2 N61P_1 (.o(UN_1_AND2_53P_I1), .i1(UN_1_AND2_59P_O), .i0(A[10]));
and2 N59P_1 (.o(UN_1_AND2_59P_O), .i1(REGSEL), .i0(SBREAD));
and2 N53P_1 (.o(UN_1_AND2_53P_O), .i1(UN_1_AND2_53P_I1), .i0(UN_1_AND2_53P_I0));
and2 N232P_1 (.o(REG32_63), .i1(UN_1_AND2_232P_I1), .i0(REGSEL));
and2 N3P_3_2 (.o(UN_3_AND2_3P_O[1]), .i1(UN_3_AND2_3P_I0[1]), .i0(UN_3_AND2_3P_I0[1]));
and2 N3P_3_1 (.i0(UN_3_AND2_3P_I0[0]), .i1(UN_3_AND2_3P_I0[0]), .o(UN_3_AND2_3P_O[0]));
and5 N90P_2 (.o(UN_2_AND5_90P_O), .i1(REG_RD_[14]), .i0(REG_WR_[9]), .i2(REG_WR_[14]), .i3(REG_RD_[15]), .i4(REG_WR_[15]));
and3 N89P_2 (.o(UN_2_AND3_89P_O), .i1(REG_WR_[7]), .i0(REG_WR_[1]), .i2(REG_WR_[8]));
and3 N70P_2 (.o(FIFO_REG), .i1(A[5]), .i0(A[4]), .i2(A[6]));
nand2 N34P_2 (.o(FIFOREG_RD_n), .i1(SBREAD), .i0(FIFOREG_REQ));
nand2 N23P_2 (.o(FIFOREG_WR_n), .i1(SBREAD_n), .i0(FIFOREG_REQ));
nand2 N15P_2 (.o(UN_2_NAND2_15P_O), .i1(A[2]), .i0(A[3]));
nand2 N5P_2 (.o(UN_2_NAND2_5P_O), .i1(A[5]), .i0(A[6]));
or2 N10P_2 (.o(UN_2_AND6_92P_I4), .i1(UN_2_OR2_10P_I1), .i0(UN_2_OR2_10P_I0));
or2 N59P_2 (.o(UN_2_OR2_58P_I1), .i1(FIFOREG_REQ), .i0(UN_2_NAND2_5P_O));
or2 N58P_2 (.o(UN_2_AND6_92P_I2), .i1(UN_2_OR2_58P_I1), .i0(UN_2_INV_6P_O));
or2 N54P_2 (.o(UN_2_AND6_92P_I0), .i1(UN_2_AND3_89P_O), .i0(REG0_31_n));
or2 N12P_2 (.o(UN_2_OR2_10P_I1), .i1(UN_2_INV_13P_O), .i0(SQCREG_REQ));
or2 N11P_2 (.o(UN_2_OR2_10P_I0), .i1(REG32_63), .i0(FIFOREG_REQ));
or2 N1P_2 (.o(UN_2_AND6_92P_I1), .i1(UN_2_AND5_90P_O), .i0(REG0_31_n));
or2 N3P_2 (.o(UN_2_AND6_92P_I3), .i1(UN_2_INV_14P_O), .i0(UN_2_NAND2_15P_O));
or2 N60P_1 (.o(UN_1_OR2_55P_I1), .i1(A[4]), .i0(A[3]));
or2 N55P_1 (.o(UN_1_AND2_53P_I0), .i1(UN_1_OR2_55P_I1), .i0(A[2]));
or2 N247P_1 (.o(REG0_15WR_n), .i1(SBREAD), .i0(REG0_31_n));
or2 N245P_1 (.o(REG0_31RD_n), .i1(SBREAD_n), .i0(REG0_31_n));
or2 N244P_1 (.o(UN_1_NOR2_283P_I0), .i1(A[8]), .i0(A[7]));
or2 N227P_1 (.o(UN_1_OR2_226P_I1), .i1(A[8]), .i0(UN_1_INV_186P_O));
or2 N226P_1 (.o(UN_1_OR2_182P_I0), .i1(UN_1_OR2_226P_I1), .i0(A[6]));
or2 N195P_1 (.o(UN_1_NOR2_283P_I1), .i1(A[10]), .i0(UN_1_INV_194P_O));
or2 N182P_1 (.o(REG0_31_n), .i1(UN_1_OR2_169P_O), .i0(UN_1_OR2_182P_I0));
or2 N169P_1 (.o(UN_1_OR2_169P_O), .i1(A[10]), .i0(A[9]));
inv N52P_2 (.o(REGSEL_n), .i(REGSEL));
inv N91P_2 (.o(DTACK_REQ_n), .i(UN_2_AND6_92P_O));
inv N68P_2 (.o(UN_2_INV_41P_I), .i(UN_2_INV_67P_O));
inv N67P_2 (.o(UN_2_INV_67P_O), .i(UN_2_INV_47P_O));
inv N51P_2 (.o(UN_2_INV_50P_I), .i(REGSEL_n));
inv N50P_2 (.o(UN_2_INV_48P_I), .i(UN_2_INV_50P_I));
inv N49P_2 (.o(UN_2_INV_47P_I), .i(UN_2_INV_48P_O));
inv N48P_2 (.o(UN_2_INV_48P_O), .i(UN_2_INV_48P_I));
inv N47P_2 (.o(UN_2_INV_47P_O), .i(UN_2_INV_47P_I));
inv N45P_2 (.o(D_REGSEL), .i(D_REGSEL_n));
inv N43P_2 (.o(D_REGSEL_n), .i(UN_2_INV_42P_O));
inv N42P_2 (.o(UN_2_INV_42P_O), .i(UN_2_INV_41P_O));
inv N41P_2 (.o(UN_2_INV_41P_O), .i(UN_2_INV_41P_I));
inv N14P_2 (.o(UN_2_INV_14P_O), .i(FIFOREG_REQ));
inv N13P_2 (.o(UN_2_INV_13P_O), .i(REG0_31_n));
inv N6P_2 (.o(UN_2_INV_6P_O), .i(REG32_63));
inv N62P_1 (.o(SBREAD), .i(SBREAD_n));
inv N348P_1 (.o(REG_WR_[4]), .i(UN_1_INV_348P_I));
inv N346P_1 (.o(REG_WR_[11]), .i(UN_1_INV_346P_I));
inv N234P_1 (.o(UN_1_INV_234P_O), .i(FIFO_REG));
inv N194P_1 (.o(UN_1_INV_194P_O), .i(A[9]));
inv N186P_1 (.o(UN_1_INV_186P_O), .i(A[7]));
inv N113P_1 (.o(CREG_REG_n), .i(UN_1_AND2_53P_O));
endmodule
`uselib

module bregs96_globals();

wire GR;
endmodule

