/* 
 *  Created:  < wittich 04/08/95>
 *  Time-stamp: <95/09/21 13:09:57 wittich>
 *  filename: /tape/snopcb/snolib_fec32/conn90/verilog_lib/verilog.v
 *  
 *  Comments: verilog model for 90 pin connector.  Simple pass-through.
 *
 *  Modification History:
 *  ------------------------------
 *  04/08/95          Created. PW.
 *  21/09/95          nuked.  back to one-sided conn 
 */

module CONN90(PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7,
    PIN8, PIN9, PIN10,PIN11, PIN12, PIN13, PIN14, PIN15, PIN16, PIN17,
    PIN18, PIN19, PIN20,PIN21, PIN22, PIN23, PIN24, PIN25, PIN26, PIN27,
    PIN28, PIN29, PIN30,PIN31, PIN32, PIN33, PIN34, PIN35, PIN36, PIN37,
    PIN38, PIN39, PIN40,PIN41, PIN42, PIN43, PIN44, PIN45, PIN46, PIN47,
    PIN48, PIN49, PIN50,PIN51, PIN52, PIN53, PIN54, PIN55, PIN56, PIN57,
    PIN58, PIN59, PIN60,PIN61, PIN62, PIN63, PIN64, PIN65, PIN66, PIN67,
    PIN68, PIN69, PIN70,PIN71, PIN72, PIN73, PIN74, PIN75, PIN76, PIN77,
    PIN78, PIN79, PIN80,PIN81, PIN82, PIN83, PIN84, PIN85, PIN86, PIN87,
 PIN88, PIN89, PIN90);

   inout PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7,
    PIN8, PIN9, PIN10;
   inout PIN11, PIN12, PIN13, PIN14, PIN15, PIN16, PIN17,
    PIN18, PIN19, PIN20;
   inout PIN21, PIN22, PIN23, PIN24, PIN25, PIN26, PIN27,
    PIN28, PIN29, PIN30;
   inout PIN31, PIN32, PIN33, PIN34, PIN35, PIN36, PIN37,
    PIN38, PIN39, PIN40;
   inout PIN41, PIN42, PIN43, PIN44, PIN45, PIN46, PIN47,
    PIN48, PIN49, PIN50;
   inout PIN51, PIN52, PIN53, PIN54, PIN55, PIN56, PIN57,
    PIN58, PIN59, PIN60;
   inout PIN61, PIN62, PIN63, PIN64, PIN65, PIN66, PIN67,
    PIN68, PIN69, PIN70;
   inout PIN71, PIN72, PIN73, PIN74, PIN75, PIN76, PIN77,
    PIN78, PIN79, PIN80;
   inout PIN81, PIN82, PIN83, PIN84, PIN85, PIN86, PIN87,
    PIN88, PIN89, PIN90;

   
   
endmodule /* CONN90 */
   


