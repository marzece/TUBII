/* 
 *  Created:  < wittich 17/08/95>
 *  Time-stamp: <95/12/06 13:58:36 wittich>
 *  filename: /tape/snopcb/snolib_fec32/mic2937a33/verilog_lib/verilog.v
 *  
 *  Comments: 5V power supply, high current.  modeled with a supply1 on
 *            output.  should I make this active only when input is high?
 *            probably not worth it.
 *
 *  Modification History:
 *  ------------------------------
 *  17/08/95          Created.
 *  06/12/95          updated for mic293blah blah blah
 */ 

module mic2937a33(INPUT, OUTPUT, GROUND);
   input INPUT,GROUND;
   output  OUTPUT;

endmodule /* mic2937a33 */

   

