/* 
 *  Created:  < wittich 14/08/95>
 *  Time-stamp: <95/08/14 14:51:50 wittich>
 *  filename: /tape/snopcb/snolib_fec32/testpoint_ls/verilog_lib/verilog.v
 *  
 *  Comments: test point dummy model.
 *
 *  Modification History:
 *  ------------------------------
 *  14/08/95          Created.
 *  12/11/95          Made sizeable.  DFC.
 * 
 */ 

module TESTPOINT_LS(A) ;
  input A;
  
endmodule /* TESTPOINT_LS */
   

