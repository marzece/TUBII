`timescale 1ns/1ns

module ports (async_delay_in, async_delay_out, async_pulse_out, caen_anpulse, caen_out, dgth, dgtl, 
    ext_ped_in, ext_ped_out, fast_anpulse, fast_comp_outh, fast_comp_outl, gtrigh_ecl, gtrigl_ecl, 
    lockout, \lockout* , \mtcd_lo* , scope_out, sync24h_ecl, sync24h_lvds, sync24l_ecl, sync24l_lvds, 
    synch_ecl, synch_lvds, syncl_ecl, syncl_lvds, sync_delay_in, sync_delay_out, sync_pulse_out, 
    tune_anpulse, tune_comp_outh, tune_comp_outl );
// generated by  HDL Direct 16.6-p001 (v16-6-112A) 9/10/2012
// on Mon Jan 19 19:23:16 2015
// from tubii_lib/PORTS/sch_1

  inout  async_delay_in;
  inout  async_delay_out;
  inout  async_pulse_out;
  inout [11:0] caen_anpulse;
  inout [7:0] caen_out;
  inout  dgth;
  inout  dgtl;
  inout  ext_ped_in;
  inout  ext_ped_out;
  inout  fast_anpulse;
  inout  fast_comp_outh;
  inout  fast_comp_outl;
  inout  gtrigh_ecl;
  inout  gtrigl_ecl;
  inout  lockout;
  inout  \lockout* ;
  inout  \mtcd_lo* ;
  inout [7:0] scope_out;
  inout  sync24h_ecl;
  inout  sync24h_lvds;
  inout  sync24l_ecl;
  inout  sync24l_lvds;
  inout  synch_ecl;
  inout  synch_lvds;
  inout  syncl_ecl;
  inout  syncl_lvds;
  inout  sync_delay_in;
  inout  sync_delay_out;
  inout  sync_pulse_out;
  inout  tune_anpulse;
  inout  tune_comp_outh;
  inout  tune_comp_outl;
  // global signal glbl.gnd;
  // global signal glbl.vtt;

  wire  unnamed_1_8merge_i149_a;
  wire  unnamed_1_8merge_i149_b;
  wire  unnamed_1_8merge_i149_c;
  wire  unnamed_1_8merge_i149_d;
  wire  unnamed_1_8merge_i149_e;
  wire  unnamed_1_8merge_i149_f;
  wire  unnamed_1_8merge_i149_g;
  wire  unnamed_1_8merge_i149_h;
  wire  unnamed_1_rsmd0805_i7_a;

  wire  gnd;
  wire  page1_gnd;
  wire [7:0] page1_scope_out;
  wire  vtt;
  wire  page1_vtt;

  assign gnd = glbl.gnd;
  assign page1_gnd = gnd;
  assign page1_scope_out[0:0] = scope_out[0:0];
  assign page1_scope_out[1:1] = scope_out[1:1];
  assign page1_scope_out[2:2] = scope_out[2:2];
  assign page1_scope_out[3:3] = scope_out[3:3];
  assign page1_scope_out[4:4] = scope_out[4:4];
  assign page1_scope_out[5:5] = scope_out[5:5];
  assign page1_scope_out[6:6] = scope_out[6:6];
  assign page1_scope_out[7:7] = scope_out[7:7];
  assign page1_scope_out[7:0] = scope_out[7:0];
  assign vtt = glbl.vtt;
  assign page1_vtt = vtt;
  assign unnamed_1_8merge_i149_a = scope_out[7:7];
  assign unnamed_1_8merge_i149_b = scope_out[6:6];
  assign unnamed_1_8merge_i149_c = scope_out[5:5];
  assign unnamed_1_8merge_i149_d = scope_out[4:4];
  assign unnamed_1_8merge_i149_e = scope_out[3:3];
  assign unnamed_1_8merge_i149_f = scope_out[2:2];
  assign unnamed_1_8merge_i149_g = scope_out[1:1];
  assign unnamed_1_8merge_i149_h = scope_out[0:0];

  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;
  assign gnd  = glbl.gnd;

// begin instances 

  rsmd0805 page1_i3  (.a({glbl.vtt}),
	.b(sync24l_ecl));

  rsmd0805 page1_i4  (.a({glbl.vtt}),
	.b(sync24h_ecl));

  ids_c10 page1_i5  (.pin1(gtrigh_ecl),
	.pin2(glbl.gnd),
	.pin3(glbl.gnd),
	.pin4(synch_ecl),
	.pin5(sync24h_ecl),
	.pin6(gtrigl_ecl),
	.pin7(glbl.gnd),
	.pin8(glbl.gnd),
	.pin9(syncl_ecl),
	.pin10(sync24l_ecl));

  rsmd0805 page1_i7  (.a(unnamed_1_rsmd0805_i7_a),
	.b(/* unconnected */));

  rsmd0805 page1_i8  (.a(unnamed_1_rsmd0805_i7_a),
	.b(/* unconnected */));

  testpoint_l page1_i24  (.a(ext_ped_out));

  testpoint_l page1_i25  (.a(glbl.gnd));

  testpoint_l page1_i26  (.a(ext_ped_in));

  testpoint_l page1_i27  (.a(glbl.gnd));

  rsmd0805 page1_i88  (.a({glbl.vtt}),
	.b(gtrigl_ecl));

  rsmd0805 page1_i89  (.a({glbl.vtt}),
	.b(gtrigh_ecl));

  testpoint_l page1_i142  (.a(unnamed_1_8merge_i149_a));

  testpoint_l page1_i143  (.a(unnamed_1_8merge_i149_b));

  testpoint_l page1_i144  (.a(unnamed_1_8merge_i149_c));

  testpoint_l page1_i145  (.a(unnamed_1_8merge_i149_d));

  testpoint_l page1_i146  (.a(unnamed_1_8merge_i149_e));

  testpoint_l page1_i147  (.a(unnamed_1_8merge_i149_g));

  testpoint_l page1_i148  (.a(unnamed_1_8merge_i149_f));

  testpoint_l page1_i150  (.a(unnamed_1_8merge_i149_h));

  translators page1_i151  ();

  caen_ports page1_i152  (.caen_anpulse(caen_anpulse[11:0]),
	.caen_out(caen_out[7:0]),
	.sync24h_lvds(sync24h_lvds),
	.sync24l_lvds(sync24l_lvds),
	.synch_lvds(synch_lvds),
	.syncl_lvds(syncl_lvds));

  comparator_ports page1_i153  (.fast_anpulse(fast_anpulse),
	.fast_comp_outh(fast_comp_outh),
	.fast_comp_outl(fast_comp_outl),
	.tune_anpulse(tune_anpulse),
	.tune_comp_outh(tune_comp_outh),
	.tune_comp_outl(tune_comp_outl));

  generic_utilities_ports page1_i154  (.async_delay_in(async_delay_in),
	.async_delay_out(async_delay_out),
	.async_pulse_out(async_pulse_out),
	.sync_delay_in(sync_delay_in),
	.sync_delay_out(sync_delay_out),
	.sync_pulse_out(sync_pulse_out));

  gt_delays_ports page1_i155  (.dgth(dgth),
	.dgtl(dgtl),
	.lockout(lockout),
	.\lockout* (\lockout* ),
	.\mtcd_lo* (\mtcd_lo* ));

  testpoint_l page1_i156  (.a(glbl.gnd));

  testpoint_l page1_i158  (.a(glbl.gnd));

  testpoint_l page1_i160  (.a(glbl.gnd));

  testpoint_l page1_i162  (.a(glbl.gnd));

  testpoint_l page1_i164  (.a(glbl.gnd));

  testpoint_l page1_i166  (.a(glbl.gnd));

  testpoint_l page1_i168  (.a(glbl.gnd));

  testpoint_l page1_i170  (.a(glbl.gnd));

endmodule // ports(sch_1) 
