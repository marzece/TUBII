// null module for a 44-pin connector 
// MSN, created 7/28/96  
// last modified:	7/29/96   


`timescale 1ns/1ns

module IDS_C34 (PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7, PIN8, PIN9, PIN10, PIN11, PIN12, PIN13, PIN14, PIN15, PIN16, PIN17, PIN18, PIN19, PIN20, PIN21, PIN22, PIN23, PIN24, PIN25, PIN26, PIN27, PIN28, PIN29, PIN30, PIN31, PIN32, PIN33, PIN34); 

        input 	PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7, PIN8, PIN9, PIN10, PIN11, PIN12, PIN13, PIN14, PIN15, PIN16, PIN17, PIN18, PIN19, PIN20, PIN21, PIN22, PIN23, PIN24, PIN25, PIN26, PIN27, PIN28, PIN29, PIN30, PIN31, PIN32, PIN33, PIN34;

endmodule

