// null module for a 14-pin connector 
// MSN, created 7/27/96  
// last modified:	7/27/96   


`timescale 1ns/1ns

module IDS_C14 (PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7, PIN8, PIN9, PIN10, PIN11, PIN12, PIN13, PIN14); 

        input 	PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7, PIN8, PIN9, PIN10, PIN11, PIN12, PIN13, PIN14;

endmodule

