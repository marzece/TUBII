/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from seq32t.xcd on Fri Oct 20 12:37:33 1995 */
/* PART 3064PQ160-100 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module sequencer32
(SDOUT, SDIN, M2, RESET_n, BXREG_WR_n, BXREG_SEL, BXREG_RD_n, BXDT, BTAG, BSEQ_RESET, BRD_STROBE, BN_ENW, BMEMREQ2_n, BMEMACK2_n, BLATCH, BFECBUSY, BDAVAIL, BCREGSEL, BCREG_REQ, BCONV_DONE, BCLKA, BCLK, BCHOLD_n, BCHIP_SEL_EN, BCAD_EN, BADC_CONVERT_n, P1, P2, P3, P6, P7, P21, P37, P38, P39, RDATA_n, RTRIG, P44, P50, P51, P70, P71, P74, P75, P76, PROGRAM_n, P81, P82, P83, P85, P94, P95, P104, P106, P107, P114, P115, P118, P119, P120, CCLK, P125, P131, P132, P133, P138, P143, P144, P151, P154, PWRDWN_n);
   output SDOUT;
   input SDIN;
   output M2;
   input RESET_n;
   input BXREG_WR_n;
   input [2:0] BXREG_SEL;
   input BXREG_RD_n;
   inout [31:0] BXDT;
   output [4:0] BTAG;
   input BSEQ_RESET;
   output BRD_STROBE;
   output [3:1] BN_ENW;
   output BMEMREQ2_n;
   input BMEMACK2_n;
   output [4:1] BLATCH;
   output BFECBUSY;
   input [32:1] BDAVAIL;
   output BCREGSEL;
   input BCREG_REQ;
   output BCONV_DONE;
   input BCLKA;
   input BCLK;
   output BCHOLD_n;
   output BCHIP_SEL_EN;
   output BCAD_EN;
   output BADC_CONVERT_n;
   inout P1;
   inout P2;
   inout P3;
   inout P6;
   inout P7;
   inout P21;
   inout P37;
   inout P38;
   inout P39;
   output RDATA_n;
   input RTRIG;
   inout P44;
   inout P50;
   inout P51;
   inout P70;
   inout P71;
   inout P74;
   inout P75;
   inout P76;
   input PROGRAM_n;
   inout P81;
   inout P82;
   inout P83;
   inout P85;
   inout P94;
   inout P95;
   inout P104;
   inout P106;
   inout P107;
   inout P114;
   inout P115;
   inout P118;
   inout P119;
   inout P120;
   input CCLK;
   inout P125;
   inout P131;
   inout P132;
   inout P133;
   inout P138;
   inout P143;
   inout P144;
   inout P151;
   inout P154;
   input PWRDWN_n;
wire [2:0] XREG_SEL;
wire [31:0] XDT;
wire [31:0] XD;
wire [4:0] TAG;
wire [32:1] LAST_SELECTED_;
wire [3:0] EO;
wire [32:1] DAVM_;
wire [32:1] DAVAIL;
wire [32:1] CS_;
wire [32:1] CHIP_MASK;
wire [32:1] CDIS;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/snolib_fec32/sequencer32/verilog_lib/sequencer32.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

fdce N115P_13_I6_1_32 (.q(CDIS[32]), .d(XD[31]), .c(N115P_13_CB), .clr(SEQ_RESET), .ce(XVDD), .gr(RESET_n));
fdce N115P_13_I6_1_31 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[30]), .q(CDIS[31]), .gr(RESET_n));
fdce N115P_13_I6_1_30 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[29]), .q(CDIS[30]), .gr(RESET_n));
fdce N115P_13_I6_1_29 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[28]), .q(CDIS[29]), .gr(RESET_n));
fdce N115P_13_I6_1_28 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[27]), .q(CDIS[28]), .gr(RESET_n));
fdce N115P_13_I6_1_27 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[26]), .q(CDIS[27]), .gr(RESET_n));
fdce N115P_13_I6_1_26 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[25]), .q(CDIS[26]), .gr(RESET_n));
fdce N115P_13_I6_1_25 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[24]), .q(CDIS[25]), .gr(RESET_n));
fdce N115P_13_I6_1_24 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[23]), .q(CDIS[24]), .gr(RESET_n));
fdce N115P_13_I6_1_23 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[22]), .q(CDIS[23]), .gr(RESET_n));
fdce N115P_13_I6_1_22 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[21]), .q(CDIS[22]), .gr(RESET_n));
fdce N115P_13_I6_1_21 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[20]), .q(CDIS[21]), .gr(RESET_n));
fdce N115P_13_I6_1_20 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[19]), .q(CDIS[20]), .gr(RESET_n));
fdce N115P_13_I6_1_19 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[18]), .q(CDIS[19]), .gr(RESET_n));
fdce N115P_13_I6_1_18 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[17]), .q(CDIS[18]), .gr(RESET_n));
fdce N115P_13_I6_1_17 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[16]), .q(CDIS[17]), .gr(RESET_n));
fdce N115P_13_I6_1_16 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[15]), .q(CDIS[16]), .gr(RESET_n));
fdce N115P_13_I6_1_15 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[14]), .q(CDIS[15]), .gr(RESET_n));
fdce N115P_13_I6_1_14 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[13]), .q(CDIS[14]), .gr(RESET_n));
fdce N115P_13_I6_1_13 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[12]), .q(CDIS[13]), .gr(RESET_n));
fdce N115P_13_I6_1_12 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[11]), .q(CDIS[12]), .gr(RESET_n));
fdce N115P_13_I6_1_11 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[10]), .q(CDIS[11]), .gr(RESET_n));
fdce N115P_13_I6_1_10 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[9]), .q(CDIS[10]), .gr(RESET_n));
fdce N115P_13_I6_1_9 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[8]), .q(CDIS[9]), .gr(RESET_n));
fdce N115P_13_I6_1_8 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[7]), .q(CDIS[8]), .gr(RESET_n));
fdce N115P_13_I6_1_7 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[6]), .q(CDIS[7]), .gr(RESET_n));
fdce N115P_13_I6_1_6 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[5]), .q(CDIS[6]), .gr(RESET_n));
fdce N115P_13_I6_1_5 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[4]), .q(CDIS[5]), .gr(RESET_n));
fdce N115P_13_I6_1_4 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[3]), .q(CDIS[4]), .gr(RESET_n));
fdce N115P_13_I6_1_3 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[2]), .q(CDIS[3]), .gr(RESET_n));
fdce N115P_13_I6_1_2 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[1]), .q(CDIS[2]), .gr(RESET_n));
fdce N115P_13_I6_1_1 (.ce(XVDD), .clr(SEQ_RESET), .c(N115P_13_CB), .d(XD[0]), .q(CDIS[1]), .gr(RESET_n));
inv N115P_13_I7_1 (.i(XREG_CDIS_WR), .o(N115P_13_CB));
and3b2 N130P_5_I30_1 (.o(N130P_5_D2), .i1(DAVM_[22]), .i0(EO[3]), .i2(DAVM_[23]));
nand2b1 N130P_5_I35_1 (.o(UN_5_X74_148_128P_I2), .i1(EO[2]), .i0(EO[3]));
and4b2 N130P_5_I34_1 (.i3(DAVM_[21]), .o(N130P_5_D5), .i1(DAVM_[20]), .i0(EO[3]), .i2(DAVM_[22]));
and4b2 N130P_5_I32_1 (.i3(DAVM_[21]), .o(N130P_5_D1), .i1(DAVM_[20]), .i0(EO[3]), .i2(DAVM_[23]));
and4b2 N130P_5_I26_1 (.i3(DAVM_[21]), .o(N130P_5_D4), .i1(DAVM_[19]), .i0(EO[3]), .i2(DAVM_[22]));
and5b1 N130P_5_I28_1 (.i4(DAVM_[21]), .i3(DAVM_[22]), .o(N130P_5_UN_1_AND5B1_I28_O), .i2(DAVM_[24]), .i0(EO[3]), .i1(DAVM_[23]));
and5b1 N130P_5_I19_1 (.i4(DAVM_[17]), .i3(DAVM_[18]), .o(N130P_5_UN_1_AND5B1_I19_O), .i2(DAVM_[20]), .i0(EO[3]), .i1(DAVM_[19]));
and5b2 N130P_5_I18_1 (.i4(DAVM_[19]), .i3(DAVM_[21]), .o(N130P_5_D0), .i1(DAVM_[18]), .i0(EO[3]), .i2(DAVM_[23]));
nor4 N130P_5_I33_1 (.i3(N130P_5_D0), .o(UN_5_NAND4_135P_I2), .i1(N130P_5_D2), .i0(N130P_5_D3), .i2(N130P_5_D1));
nor4 N130P_5_I16_1 (.i3(N130P_5_D8), .o(UN_5_NAND4_137P_I0), .i1(N130P_5_D10), .i0(N130P_5_D11), .i2(N130P_5_D9));
nor4 N130P_5_I15_1 (.i3(N130P_5_D4), .o(UN_5_NAND4_136P_I2), .i1(N130P_5_D6), .i0(N130P_5_D7), .i2(N130P_5_D5));
nand2 N130P_5_I20_1 (.o(EO[2]), .i1(N130P_5_UN_1_AND5B1_I19_O), .i0(N130P_5_UN_1_AND5B1_I28_O));
nor2 N130P_5_I29_1 (.o(N130P_5_D11), .i1(DAVM_[24]), .i0(EO[3]));
nor2 N130P_5_I27_1 (.o(N130P_5_D7), .i1(DAVM_[24]), .i0(EO[3]));
nor2 N130P_5_I24_1 (.o(N130P_5_D9), .i1(DAVM_[22]), .i0(EO[3]));
nor2 N130P_5_I25_1 (.o(N130P_5_D6), .i1(DAVM_[23]), .i0(EO[3]));
nor2 N130P_5_I23_1 (.o(N130P_5_D3), .i1(DAVM_[24]), .i0(EO[3]));
nor2 N130P_5_I21_1 (.o(N130P_5_D10), .i1(DAVM_[23]), .i0(EO[3]));
nor2 N130P_5_I17_1 (.o(N130P_5_D8), .i1(DAVM_[21]), .i0(EO[3]));
and3b2 N129P_5_I30_1 (.o(N129P_5_D2), .i1(DAVM_[6]), .i0(EO[1]), .i2(DAVM_[7]));
nand2b1 N129P_5_I35_1 (.o(UN_5_X74_148_128P_I0), .i1(EO[0]), .i0(EO[1]));
and4b2 N129P_5_I34_1 (.i3(DAVM_[5]), .o(N129P_5_D5), .i1(DAVM_[4]), .i0(EO[1]), .i2(DAVM_[6]));
and4b2 N129P_5_I32_1 (.i3(DAVM_[5]), .o(N129P_5_D1), .i1(DAVM_[4]), .i0(EO[1]), .i2(DAVM_[7]));
and4b2 N129P_5_I26_1 (.i3(DAVM_[5]), .o(N129P_5_D4), .i1(DAVM_[3]), .i0(EO[1]), .i2(DAVM_[6]));
and5b1 N129P_5_I28_1 (.i4(DAVM_[5]), .i3(DAVM_[6]), .o(N129P_5_UN_1_AND5B1_I28_O), .i2(DAVM_[8]), .i0(EO[1]), .i1(DAVM_[7]));
and5b1 N129P_5_I19_1 (.i4(DAVM_[1]), .i3(DAVM_[2]), .o(N129P_5_UN_1_AND5B1_I19_O), .i2(DAVM_[4]), .i0(EO[1]), .i1(DAVM_[3]));
and5b2 N129P_5_I18_1 (.i4(DAVM_[3]), .i3(DAVM_[5]), .o(N129P_5_D0), .i1(DAVM_[2]), .i0(EO[1]), .i2(DAVM_[7]));
nor4 N129P_5_I33_1 (.i3(N129P_5_D0), .o(UN_5_NAND4_135P_I0), .i1(N129P_5_D2), .i0(N129P_5_D3), .i2(N129P_5_D1));
nor4 N129P_5_I16_1 (.i3(N129P_5_D8), .o(UN_5_NAND4_137P_I1), .i1(N129P_5_D10), .i0(N129P_5_D11), .i2(N129P_5_D9));
nor4 N129P_5_I15_1 (.i3(N129P_5_D4), .o(UN_5_NAND4_136P_I1), .i1(N129P_5_D6), .i0(N129P_5_D7), .i2(N129P_5_D5));
nand2 N129P_5_I20_1 (.o(EO[0]), .i1(N129P_5_UN_1_AND5B1_I19_O), .i0(N129P_5_UN_1_AND5B1_I28_O));
nor2 N129P_5_I29_1 (.o(N129P_5_D11), .i1(DAVM_[8]), .i0(EO[1]));
nor2 N129P_5_I27_1 (.o(N129P_5_D7), .i1(DAVM_[8]), .i0(EO[1]));
nor2 N129P_5_I24_1 (.o(N129P_5_D9), .i1(DAVM_[6]), .i0(EO[1]));
nor2 N129P_5_I25_1 (.o(N129P_5_D6), .i1(DAVM_[7]), .i0(EO[1]));
nor2 N129P_5_I23_1 (.o(N129P_5_D3), .i1(DAVM_[8]), .i0(EO[1]));
nor2 N129P_5_I21_1 (.o(N129P_5_D10), .i1(DAVM_[7]), .i0(EO[1]));
nor2 N129P_5_I17_1 (.o(N129P_5_D8), .i1(DAVM_[5]), .i0(EO[1]));
and3b2 N131P_5_I30_1 (.o(N131P_5_D2), .i1(DAVM_[14]), .i0(EO[2]), .i2(DAVM_[15]));
nand2b1 N131P_5_I35_1 (.o(UN_5_X74_148_128P_I1), .i1(EO[1]), .i0(EO[2]));
and4b2 N131P_5_I34_1 (.i3(DAVM_[13]), .o(N131P_5_D5), .i1(DAVM_[12]), .i0(EO[2]), .i2(DAVM_[14]));
and4b2 N131P_5_I32_1 (.i3(DAVM_[13]), .o(N131P_5_D1), .i1(DAVM_[12]), .i0(EO[2]), .i2(DAVM_[15]));
and4b2 N131P_5_I26_1 (.i3(DAVM_[13]), .o(N131P_5_D4), .i1(DAVM_[11]), .i0(EO[2]), .i2(DAVM_[14]));
and5b1 N131P_5_I28_1 (.i4(DAVM_[13]), .i3(DAVM_[14]), .o(N131P_5_UN_1_AND5B1_I28_O), .i2(DAVM_[16]), .i0(EO[2]), .i1(DAVM_[15]));
and5b1 N131P_5_I19_1 (.i4(DAVM_[9]), .i3(DAVM_[10]), .o(N131P_5_UN_1_AND5B1_I19_O), .i2(DAVM_[12]), .i0(EO[2]), .i1(DAVM_[11]));
and5b2 N131P_5_I18_1 (.i4(DAVM_[11]), .i3(DAVM_[13]), .o(N131P_5_D0), .i1(DAVM_[10]), .i0(EO[2]), .i2(DAVM_[15]));
nor4 N131P_5_I33_1 (.i3(N131P_5_D0), .o(UN_5_NAND4_135P_I1), .i1(N131P_5_D2), .i0(N131P_5_D3), .i2(N131P_5_D1));
nor4 N131P_5_I16_1 (.i3(N131P_5_D8), .o(UN_5_NAND4_137P_I2), .i1(N131P_5_D10), .i0(N131P_5_D11), .i2(N131P_5_D9));
nor4 N131P_5_I15_1 (.i3(N131P_5_D4), .o(UN_5_NAND4_136P_I0), .i1(N131P_5_D6), .i0(N131P_5_D7), .i2(N131P_5_D5));
nand2 N131P_5_I20_1 (.o(EO[1]), .i1(N131P_5_UN_1_AND5B1_I19_O), .i0(N131P_5_UN_1_AND5B1_I28_O));
nor2 N131P_5_I29_1 (.o(N131P_5_D11), .i1(DAVM_[16]), .i0(EO[2]));
nor2 N131P_5_I27_1 (.o(N131P_5_D7), .i1(DAVM_[16]), .i0(EO[2]));
nor2 N131P_5_I24_1 (.o(N131P_5_D9), .i1(DAVM_[14]), .i0(EO[2]));
nor2 N131P_5_I25_1 (.o(N131P_5_D6), .i1(DAVM_[15]), .i0(EO[2]));
nor2 N131P_5_I23_1 (.o(N131P_5_D3), .i1(DAVM_[16]), .i0(EO[2]));
nor2 N131P_5_I21_1 (.o(N131P_5_D10), .i1(DAVM_[15]), .i0(EO[2]));
nor2 N131P_5_I17_1 (.o(N131P_5_D8), .i1(DAVM_[13]), .i0(EO[2]));
and3b2 N128P_5_I30_1 (.o(N128P_5_D2), .i1(XVDD), .i0(XGND), .i2(XVDD));
nand2b1 N128P_5_I35_1 (.o(N128P_5_GS), .i1(N128P_5_EO), .i0(XGND));
and4b2 N128P_5_I34_1 (.i3(XVDD), .o(N128P_5_D5), .i1(UN_5_X74_148_127P_GS), .i0(XGND), .i2(XVDD));
and4b2 N128P_5_I32_1 (.i3(XVDD), .o(N128P_5_D1), .i1(UN_5_X74_148_127P_GS), .i0(XGND), .i2(XVDD));
and4b2 N128P_5_I26_1 (.i3(XVDD), .o(N128P_5_D4), .i1(UN_5_X74_148_128P_I2), .i0(XGND), .i2(XVDD));
and5b1 N128P_5_I28_1 (.i4(XVDD), .i3(XVDD), .o(N128P_5_UN_1_AND5B1_I28_O), .i2(XVDD), .i0(XGND), .i1(XVDD));
and5b1 N128P_5_I19_1 (.i4(UN_5_X74_148_128P_I0), .i3(UN_5_X74_148_128P_I1), .o(N128P_5_UN_1_AND5B1_I19_O), .i2(UN_5_X74_148_127P_GS), .i0(XGND), .i1(UN_5_X74_148_128P_I2));
and5b2 N128P_5_I18_1 (.i4(UN_5_X74_148_128P_I2), .i3(XVDD), .o(N128P_5_D0), .i1(UN_5_X74_148_128P_I1), .i0(XGND), .i2(XVDD));
nor4 N128P_5_I33_1 (.i3(N128P_5_D0), .o(UN_5_INV_149P_I), .i1(N128P_5_D2), .i0(N128P_5_D3), .i2(N128P_5_D1));
nor4 N128P_5_I16_1 (.i3(N128P_5_D8), .o(N128P_5_A2), .i1(N128P_5_D10), .i0(N128P_5_D11), .i2(N128P_5_D9));
nor4 N128P_5_I15_1 (.i3(N128P_5_D4), .o(UN_5_INV_148P_I), .i1(N128P_5_D6), .i0(N128P_5_D7), .i2(N128P_5_D5));
nand2 N128P_5_I20_1 (.o(N128P_5_EO), .i1(N128P_5_UN_1_AND5B1_I19_O), .i0(N128P_5_UN_1_AND5B1_I28_O));
nor2 N128P_5_I29_1 (.o(N128P_5_D11), .i1(XVDD), .i0(XGND));
nor2 N128P_5_I27_1 (.o(N128P_5_D7), .i1(XVDD), .i0(XGND));
nor2 N128P_5_I24_1 (.o(N128P_5_D9), .i1(XVDD), .i0(XGND));
nor2 N128P_5_I25_1 (.o(N128P_5_D6), .i1(XVDD), .i0(XGND));
nor2 N128P_5_I23_1 (.o(N128P_5_D3), .i1(XVDD), .i0(XGND));
nor2 N128P_5_I21_1 (.o(N128P_5_D10), .i1(XVDD), .i0(XGND));
nor2 N128P_5_I17_1 (.o(N128P_5_D8), .i1(XVDD), .i0(XGND));
and3b2 N127P_5_I30_1 (.o(N127P_5_D2), .i1(DAVM_[30]), .i0(XGND), .i2(DAVM_[31]));
nand2b1 N127P_5_I35_1 (.o(UN_5_X74_148_127P_GS), .i1(EO[3]), .i0(XGND));
and4b2 N127P_5_I34_1 (.i3(DAVM_[29]), .o(N127P_5_D5), .i1(DAVM_[28]), .i0(XGND), .i2(DAVM_[30]));
and4b2 N127P_5_I32_1 (.i3(DAVM_[29]), .o(N127P_5_D1), .i1(DAVM_[28]), .i0(XGND), .i2(DAVM_[31]));
and4b2 N127P_5_I26_1 (.i3(DAVM_[29]), .o(N127P_5_D4), .i1(DAVM_[27]), .i0(XGND), .i2(DAVM_[30]));
and5b1 N127P_5_I28_1 (.i4(DAVM_[29]), .i3(DAVM_[30]), .o(N127P_5_UN_1_AND5B1_I28_O), .i2(DAVM_[32]), .i0(XGND), .i1(DAVM_[31]));
and5b1 N127P_5_I19_1 (.i4(DAVM_[25]), .i3(DAVM_[26]), .o(N127P_5_UN_1_AND5B1_I19_O), .i2(DAVM_[28]), .i0(XGND), .i1(DAVM_[27]));
and5b2 N127P_5_I18_1 (.i4(DAVM_[27]), .i3(DAVM_[29]), .o(N127P_5_D0), .i1(DAVM_[26]), .i0(XGND), .i2(DAVM_[31]));
nor4 N127P_5_I33_1 (.i3(N127P_5_D0), .o(UN_5_NAND4_135P_I3), .i1(N127P_5_D2), .i0(N127P_5_D3), .i2(N127P_5_D1));
nor4 N127P_5_I16_1 (.i3(N127P_5_D8), .o(UN_5_NAND4_137P_I3), .i1(N127P_5_D10), .i0(N127P_5_D11), .i2(N127P_5_D9));
nor4 N127P_5_I15_1 (.i3(N127P_5_D4), .o(UN_5_NAND4_136P_I3), .i1(N127P_5_D6), .i0(N127P_5_D7), .i2(N127P_5_D5));
nand2 N127P_5_I20_1 (.o(EO[3]), .i1(N127P_5_UN_1_AND5B1_I19_O), .i0(N127P_5_UN_1_AND5B1_I28_O));
nor2 N127P_5_I29_1 (.o(N127P_5_D11), .i1(DAVM_[32]), .i0(XGND));
nor2 N127P_5_I27_1 (.o(N127P_5_D7), .i1(DAVM_[32]), .i0(XGND));
nor2 N127P_5_I24_1 (.o(N127P_5_D9), .i1(DAVM_[30]), .i0(XGND));
nor2 N127P_5_I25_1 (.o(N127P_5_D6), .i1(DAVM_[31]), .i0(XGND));
nor2 N127P_5_I23_1 (.o(N127P_5_D3), .i1(DAVM_[32]), .i0(XGND));
nor2 N127P_5_I21_1 (.o(N127P_5_D10), .i1(DAVM_[31]), .i0(XGND));
nor2 N127P_5_I17_1 (.o(N127P_5_D8), .i1(DAVM_[29]), .i0(XGND));
and3b2 N29P_13_I16_1 (.o(N29P_13_E), .i1(XREG_RD_n), .i0(XGND), .i2(XVDD));
nand4b1 N29P_13_I22_1 (.i3(N29P_13_E), .o(N29P_13_Y5), .i2(XREG_SEL[2]), .i0(XREG_SEL[1]), .i1(XREG_SEL[0]));
nand4b1 N29P_13_I18_1 (.i3(N29P_13_E), .o(N29P_13_Y3), .i2(XREG_SEL[0]), .i0(XREG_SEL[2]), .i1(XREG_SEL[1]));
nand4b1 N29P_13_I15_1 (.i3(N29P_13_E), .o(N29P_13_Y6), .i2(XREG_SEL[2]), .i0(XREG_SEL[0]), .i1(XREG_SEL[1]));
nand4b3 N29P_13_I23_1 (.i3(N29P_13_E), .o(XREG_INCS_RD_n), .i2(XREG_SEL[1]), .i1(XREG_SEL[2]), .i0(XREG_SEL[0]));
nand4b2 N29P_13_I25_1 (.i3(N29P_13_E), .o(XREG_DAV_RD_n), .i1(XREG_SEL[0]), .i0(XREG_SEL[2]), .i2(XREG_SEL[1]));
nand4b2 N29P_13_I21_1 (.i3(N29P_13_E), .o(XREG_OUTCS_RD_n), .i1(XREG_SEL[1]), .i0(XREG_SEL[2]), .i2(XREG_SEL[0]));
nand4b2 N29P_13_I20_1 (.i3(N29P_13_E), .o(N29P_13_Y4), .i1(XREG_SEL[0]), .i0(XREG_SEL[1]), .i2(XREG_SEL[2]));
nand4 N29P_13_I17_1 (.i3(N29P_13_E), .o(N29P_13_Y7), .i1(XREG_SEL[1]), .i0(XREG_SEL[2]), .i2(XREG_SEL[0]));
and3b2 N28P_13_I16_1 (.o(N28P_13_E), .i1(XREG_WR_n), .i0(XGND), .i2(XVDD));
nand4b1 N28P_13_I22_1 (.i3(N28P_13_E), .o(N28P_13_Y5), .i2(XREG_SEL[2]), .i0(XREG_SEL[1]), .i1(XREG_SEL[0]));
nand4b1 N28P_13_I18_1 (.i3(N28P_13_E), .o(N28P_13_Y3), .i2(XREG_SEL[0]), .i0(XREG_SEL[2]), .i1(XREG_SEL[1]));
nand4b1 N28P_13_I15_1 (.i3(N28P_13_E), .o(N28P_13_Y6), .i2(XREG_SEL[2]), .i0(XREG_SEL[0]), .i1(XREG_SEL[1]));
nand4b3 N28P_13_I23_1 (.i3(N28P_13_E), .o(N28P_13_Y0), .i2(XREG_SEL[1]), .i1(XREG_SEL[2]), .i0(XREG_SEL[0]));
nand4b2 N28P_13_I25_1 (.i3(N28P_13_E), .o(N28P_13_Y2), .i1(XREG_SEL[0]), .i0(XREG_SEL[2]), .i2(XREG_SEL[1]));
nand4b2 N28P_13_I21_1 (.i3(N28P_13_E), .o(N28P_13_Y1), .i1(XREG_SEL[1]), .i0(XREG_SEL[2]), .i2(XREG_SEL[0]));
nand4b2 N28P_13_I20_1 (.i3(N28P_13_E), .o(UN_13_ACLK_110P_I), .i1(XREG_SEL[0]), .i0(XREG_SEL[1]), .i2(XREG_SEL[2]));
nand4 N28P_13_I17_1 (.i3(N28P_13_E), .o(N28P_13_Y7), .i1(XREG_SEL[1]), .i0(XREG_SEL[2]), .i2(XREG_SEL[0]));
and3b2 N43P_4_I16_1 (.o(N43P_4_E), .i1(TAG[4]), .i0(TAG[3]), .i2(CHIP_SEL_EN));
nand4b1 N43P_4_I22_1 (.i3(N43P_4_E), .o(CS_[6]), .i2(TAG[2]), .i0(TAG[1]), .i1(TAG[0]));
nand4b1 N43P_4_I18_1 (.i3(N43P_4_E), .o(CS_[4]), .i2(TAG[0]), .i0(TAG[2]), .i1(TAG[1]));
nand4b1 N43P_4_I15_1 (.i3(N43P_4_E), .o(CS_[7]), .i2(TAG[2]), .i0(TAG[0]), .i1(TAG[1]));
nand4b3 N43P_4_I23_1 (.i3(N43P_4_E), .o(CS_[1]), .i2(TAG[1]), .i1(TAG[2]), .i0(TAG[0]));
nand4b2 N43P_4_I25_1 (.i3(N43P_4_E), .o(CS_[3]), .i1(TAG[0]), .i0(TAG[2]), .i2(TAG[1]));
nand4b2 N43P_4_I21_1 (.i3(N43P_4_E), .o(CS_[2]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
nand4b2 N43P_4_I20_1 (.i3(N43P_4_E), .o(CS_[5]), .i1(TAG[0]), .i0(TAG[1]), .i2(TAG[2]));
nand4 N43P_4_I17_1 (.i3(N43P_4_E), .o(CS_[8]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
and3b2 N6P_4_I16_1 (.o(N6P_4_E), .i1(UN_4_INV_77P_O), .i0(UN_4_INV_76P_O), .i2(CHIP_SEL_EN));
nand4b1 N6P_4_I22_1 (.i3(N6P_4_E), .o(CS_[30]), .i2(TAG[2]), .i0(TAG[1]), .i1(TAG[0]));
nand4b1 N6P_4_I18_1 (.i3(N6P_4_E), .o(CS_[28]), .i2(TAG[0]), .i0(TAG[2]), .i1(TAG[1]));
nand4b1 N6P_4_I15_1 (.i3(N6P_4_E), .o(CS_[31]), .i2(TAG[2]), .i0(TAG[0]), .i1(TAG[1]));
nand4b3 N6P_4_I23_1 (.i3(N6P_4_E), .o(CS_[25]), .i2(TAG[1]), .i1(TAG[2]), .i0(TAG[0]));
nand4b2 N6P_4_I25_1 (.i3(N6P_4_E), .o(CS_[27]), .i1(TAG[0]), .i0(TAG[2]), .i2(TAG[1]));
nand4b2 N6P_4_I21_1 (.i3(N6P_4_E), .o(CS_[26]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
nand4b2 N6P_4_I20_1 (.i3(N6P_4_E), .o(CS_[29]), .i1(TAG[0]), .i0(TAG[1]), .i2(TAG[2]));
nand4 N6P_4_I17_1 (.i3(N6P_4_E), .o(CS_[32]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
and3b2 N7P_4_I16_1 (.o(N7P_4_E), .i1(UN_4_INV_77P_O), .i0(TAG[3]), .i2(CHIP_SEL_EN));
nand4b1 N7P_4_I22_1 (.i3(N7P_4_E), .o(CS_[22]), .i2(TAG[2]), .i0(TAG[1]), .i1(TAG[0]));
nand4b1 N7P_4_I18_1 (.i3(N7P_4_E), .o(CS_[20]), .i2(TAG[0]), .i0(TAG[2]), .i1(TAG[1]));
nand4b1 N7P_4_I15_1 (.i3(N7P_4_E), .o(CS_[23]), .i2(TAG[2]), .i0(TAG[0]), .i1(TAG[1]));
nand4b3 N7P_4_I23_1 (.i3(N7P_4_E), .o(CS_[17]), .i2(TAG[1]), .i1(TAG[2]), .i0(TAG[0]));
nand4b2 N7P_4_I25_1 (.i3(N7P_4_E), .o(CS_[19]), .i1(TAG[0]), .i0(TAG[2]), .i2(TAG[1]));
nand4b2 N7P_4_I21_1 (.i3(N7P_4_E), .o(CS_[18]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
nand4b2 N7P_4_I20_1 (.i3(N7P_4_E), .o(CS_[21]), .i1(TAG[0]), .i0(TAG[1]), .i2(TAG[2]));
nand4 N7P_4_I17_1 (.i3(N7P_4_E), .o(CS_[24]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
and3b2 N8P_4_I16_1 (.o(N8P_4_E), .i1(UN_4_INV_76P_O), .i0(TAG[4]), .i2(CHIP_SEL_EN));
nand4b1 N8P_4_I22_1 (.i3(N8P_4_E), .o(CS_[14]), .i2(TAG[2]), .i0(TAG[1]), .i1(TAG[0]));
nand4b1 N8P_4_I18_1 (.i3(N8P_4_E), .o(CS_[12]), .i2(TAG[0]), .i0(TAG[2]), .i1(TAG[1]));
nand4b1 N8P_4_I15_1 (.i3(N8P_4_E), .o(CS_[15]), .i2(TAG[2]), .i0(TAG[0]), .i1(TAG[1]));
nand4b3 N8P_4_I23_1 (.i3(N8P_4_E), .o(CS_[9]), .i2(TAG[1]), .i1(TAG[2]), .i0(TAG[0]));
nand4b2 N8P_4_I25_1 (.i3(N8P_4_E), .o(CS_[11]), .i1(TAG[0]), .i0(TAG[2]), .i2(TAG[1]));
nand4b2 N8P_4_I21_1 (.i3(N8P_4_E), .o(CS_[10]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
nand4b2 N8P_4_I20_1 (.i3(N8P_4_E), .o(CS_[13]), .i1(TAG[0]), .i0(TAG[1]), .i2(TAG[2]));
nand4 N8P_4_I17_1 (.i3(N8P_4_E), .o(CS_[16]), .i1(TAG[1]), .i0(TAG[2]), .i2(TAG[0]));
fdce N99P_8_I8_1 (.q(LAST_SELECTED_[21]), .d(DAVAIL[21]), .c(CS_[21]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N89P_8_I8_1 (.q(LAST_SELECTED_[8]), .d(DAVAIL[8]), .c(CS_[8]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N86P_8_I8_1 (.q(LAST_SELECTED_[9]), .d(DAVAIL[9]), .c(CS_[9]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N83P_8_I8_1 (.q(LAST_SELECTED_[10]), .d(DAVAIL[10]), .c(CS_[10]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N80P_8_I8_1 (.q(LAST_SELECTED_[11]), .d(DAVAIL[11]), .c(CS_[11]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N74P_8_I8_1 (.q(LAST_SELECTED_[13]), .d(DAVAIL[13]), .c(CS_[13]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N71P_8_I8_1 (.q(LAST_SELECTED_[14]), .d(DAVAIL[14]), .c(CS_[14]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N178P_8_I8_1 (.q(LAST_SELECTED_[2]), .d(DAVAIL[2]), .c(CS_[2]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N163P_8_I8_1 (.q(LAST_SELECTED_[28]), .d(DAVAIL[28]), .c(CS_[28]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N160P_8_I8_1 (.q(LAST_SELECTED_[29]), .d(DAVAIL[29]), .c(CS_[29]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N154P_8_I8_1 (.q(LAST_SELECTED_[31]), .d(DAVAIL[31]), .c(CS_[31]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N151P_8_I8_1 (.q(LAST_SELECTED_[32]), .d(DAVAIL[32]), .c(CS_[32]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N117P_8_I8_1 (.q(LAST_SELECTED_[15]), .d(DAVAIL[15]), .c(CS_[15]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N114P_8_I8_1 (.q(LAST_SELECTED_[16]), .d(DAVAIL[16]), .c(CS_[16]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N111P_8_I8_1 (.q(LAST_SELECTED_[17]), .d(DAVAIL[17]), .c(CS_[17]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N108P_8_I8_1 (.q(LAST_SELECTED_[18]), .d(DAVAIL[18]), .c(CS_[18]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N105P_8_I8_1 (.q(LAST_SELECTED_[19]), .d(DAVAIL[19]), .c(CS_[19]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N102P_8_I8_1 (.q(LAST_SELECTED_[20]), .d(DAVAIL[20]), .c(CS_[20]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N130P_8_I8_1 (.q(LAST_SELECTED_[26]), .d(DAVAIL[26]), .c(CS_[26]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N77P_8_I8_1 (.q(LAST_SELECTED_[12]), .d(DAVAIL[12]), .c(CS_[12]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N181P_8_I8_1 (.q(LAST_SELECTED_[3]), .d(DAVAIL[3]), .c(CS_[3]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N176P_8_I8_1 (.q(LAST_SELECTED_[1]), .d(DAVAIL[1]), .c(CS_[1]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N193P_8_I8_1 (.q(LAST_SELECTED_[7]), .d(DAVAIL[7]), .c(CS_[7]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N190P_8_I8_1 (.q(LAST_SELECTED_[6]), .d(DAVAIL[6]), .c(CS_[6]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N187P_8_I8_1 (.q(LAST_SELECTED_[5]), .d(DAVAIL[5]), .c(CS_[5]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N184P_8_I8_1 (.q(LAST_SELECTED_[4]), .d(DAVAIL[4]), .c(CS_[4]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N157P_8_I8_1 (.q(LAST_SELECTED_[30]), .d(DAVAIL[30]), .c(CS_[30]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N142P_8_I8_1 (.q(LAST_SELECTED_[22]), .d(DAVAIL[22]), .c(CS_[22]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N139P_8_I8_1 (.q(LAST_SELECTED_[23]), .d(DAVAIL[23]), .c(CS_[23]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N136P_8_I8_1 (.q(LAST_SELECTED_[24]), .d(DAVAIL[24]), .c(CS_[24]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N133P_8_I8_1 (.q(LAST_SELECTED_[25]), .d(DAVAIL[25]), .c(CS_[25]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N127P_8_I8_1 (.q(LAST_SELECTED_[27]), .d(DAVAIL[27]), .c(CS_[27]), .clr(DAV_n), .ce(XVDD), .gr(RESET_n));
fdce N170P_3_I8_1 (.q(UN_3_FDC_164P_D), .d(CAD_EN), .c(CLK), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N166P_3_I8_1 (.q(UN_3_FDC_166P_Q), .d(UN_3_FDC_165P_Q), .c(CLK), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N165P_3_I8_1 (.q(UN_3_FDC_165P_Q), .d(UN_3_FDC_164P_Q), .c(CLK), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N164P_3_I8_1 (.q(UN_3_FDC_164P_Q), .d(UN_3_FDC_164P_D), .c(CLK), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N144P_3_I8_1 (.q(UN_3_FDC_144P_Q), .d(UN_3_FDC_142P_C), .c(CLK), .clr(SEQ_RESET), .ce(XVDD), .gr(RESET_n));
fdce N142P_3_I8_1 (.q(UN_3_FDC_142P_Q), .d(UN_3_FDC_142P_D), .c(UN_3_FDC_142P_C), .clr(UN_3_FDC_142P_CLR), .ce(XVDD), .gr(RESET_n));
fdce N139P_3_I8_1 (.q(UN_3_FDC_139P_Q), .d(UN_3_FDC_128P_C), .c(UN_3_FDC_142P_D), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N136P_3_I8_1 (.q(UN_3_FDC_136P_Q), .d(UN_3_FDC_133P_C), .c(UN_3_FDC_136P_C), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N133P_3_I8_1 (.q(UN_3_FDC_133P_Q), .d(UN_3_FDC_133P_D), .c(UN_3_FDC_133P_C), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N132P_3_I8_1 (.q(UN_3_FDC_131P_D), .d(UN_3_FDC_133P_Q), .c(CLK), .clr(UN_3_FDC_132P_CLR), .ce(XVDD), .gr(RESET_n));
fdce N131P_3_I8_1 (.q(UN_3_FDC_131P_Q), .d(UN_3_FDC_131P_D), .c(CLK), .clr(SEQ_RESET), .ce(XVDD), .gr(RESET_n));
fdce N128P_3_I8_1 (.q(UN_3_FDC_128P_Q), .d(UN_3_FDC_136P_C), .c(UN_3_FDC_128P_C), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N127P_3_I8_1 (.q(UN_3_FDC_127P_Q), .d(ADC_CONVERT), .c(UN_3_FDC_128P_C), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N126P_3_I8_1 (.q(ADC_CONVERT), .d(UN_3_FDC_126P_D), .c(UN_3_FDC_128P_C), .clr(CONV_DONE), .ce(XVDD), .gr(RESET_n));
fdce N179P_2_I8_1 (.q(UN_2_AND3_209P_I2), .d(UN_2_AND3_208P_I1), .c(UN_2_FDC_171P_C), .clr(MEMCLR_n), .ce(XVDD), .gr(RESET_n));
fdce N172P_2_I8_1 (.q(UN_2_AND2_210P_I1), .d(UN_2_AND3_209P_I2), .c(UN_2_FDC_171P_C), .clr(MEMCLR_n), .ce(XVDD), .gr(RESET_n));
fdce N171P_2_I8_1 (.q(UN_2_FDC_171P_Q), .d(UN_2_AND2_210P_I1), .c(UN_2_FDC_171P_C), .clr(MEMCLR_n), .ce(XVDD), .gr(RESET_n));
fdce N180P_2_I8_1 (.q(UN_2_AND3_208P_I1), .d(UN_2_FDC_180P_D), .c(LATCH3), .clr(MEMCLR_n), .ce(XVDD), .gr(RESET_n));
fdce N213P_1_I8_1 (.q(UN_1_FDC_213P_Q), .d(CHIP_SEL_EN), .c(CLK), .clr(UN_1_AND2_262P_O), .ce(XVDD), .gr(RESET_n));
fdce N205P_1_I8_1 (.q(UN_1_FDC_205P_Q), .d(SEQ_RESET_n), .c(CREG_REQ), .clr(UN_1_FDC_205P_CLR), .ce(XVDD), .gr(RESET_n));
fdce N203P_1_I8_1 (.q(CAD_EN), .d(UPSTART), .c(CLK), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N202P_1_I8_1 (.q(CHIP_SEL_EN), .d(CAD_EN), .c(CLK_n), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N201P_1_I8_1 (.q(LATCH1), .d(CHIP_SEL_EN), .c(RD_STROBE), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N200P_1_I8_1 (.q(LATCH2), .d(LATCH1), .c(RD_STROBE), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N199P_1_I8_1 (.q(LATCH3), .d(LATCH2), .c(RD_STROBE), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N198P_1_I8_1 (.q(LATCH4), .d(LATCH3), .c(RD_STROBE), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N192P_1_I8_1 (.q(FECSTART), .d(UN_1_FDC_192P_D), .c(CLK), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N191P_1_I8_1 (.q(FECSEL_n), .d(UN_1_FDC_191P_D), .c(CLK), .clr(CDONE), .ce(XVDD), .gr(RESET_n));
fdce N183P_1_I8_1 (.q(UN_1_FDC_183P_Q), .d(UN_1_FDC_183P_D), .c(CLK), .clr(UN_1_FDC_183P_CLR), .ce(XVDD), .gr(RESET_n));
pullup1 N121P_13_32 (.o(XDT[31]));
pullup1 N121P_13_31 (.o(XDT[30]));
pullup1 N121P_13_30 (.o(XDT[29]));
pullup1 N121P_13_29 (.o(XDT[28]));
pullup1 N121P_13_28 (.o(XDT[27]));
pullup1 N121P_13_27 (.o(XDT[26]));
pullup1 N121P_13_26 (.o(XDT[25]));
pullup1 N121P_13_25 (.o(XDT[24]));
pullup1 N121P_13_24 (.o(XDT[23]));
pullup1 N121P_13_23 (.o(XDT[22]));
pullup1 N121P_13_22 (.o(XDT[21]));
pullup1 N121P_13_21 (.o(XDT[20]));
pullup1 N121P_13_20 (.o(XDT[19]));
pullup1 N121P_13_19 (.o(XDT[18]));
pullup1 N121P_13_18 (.o(XDT[17]));
pullup1 N121P_13_17 (.o(XDT[16]));
pullup1 N121P_13_16 (.o(XDT[15]));
pullup1 N121P_13_15 (.o(XDT[14]));
pullup1 N121P_13_14 (.o(XDT[13]));
pullup1 N121P_13_13 (.o(XDT[12]));
pullup1 N121P_13_12 (.o(XDT[11]));
pullup1 N121P_13_11 (.o(XDT[10]));
pullup1 N121P_13_10 (.o(XDT[9]));
pullup1 N121P_13_9 (.o(XDT[8]));
pullup1 N121P_13_8 (.o(XDT[7]));
pullup1 N121P_13_7 (.o(XDT[6]));
pullup1 N121P_13_6 (.o(XDT[5]));
pullup1 N121P_13_5 (.o(XDT[4]));
pullup1 N121P_13_4 (.o(XDT[3]));
pullup1 N121P_13_3 (.o(XDT[2]));
pullup1 N121P_13_2 (.o(XDT[1]));
pullup1 N121P_13_1 (.o(XDT[0]));
buft N94P_13_8 (.i(CHOLD_n), .o(XDT[15]), .t(XREG_OUTCS_RD_n));
buft N94P_13_7 (.t(XREG_OUTCS_RD_n), .o(XDT[14]), .i(ENW3_n));
buft N94P_13_6 (.t(XREG_OUTCS_RD_n), .o(XDT[13]), .i(ENW2_n));
buft N94P_13_5 (.t(XREG_OUTCS_RD_n), .o(XDT[12]), .i(ENW1_n));
buft N94P_13_4 (.t(XREG_OUTCS_RD_n), .o(XDT[11]), .i(MEMREQ2_n));
buft N94P_13_3 (.t(XREG_OUTCS_RD_n), .o(XDT[10]), .i(CAD_EN));
buft N94P_13_2 (.t(XREG_OUTCS_RD_n), .o(XDT[9]), .i(ADC_CONVERT_n));
buft N94P_13_1 (.t(XREG_OUTCS_RD_n), .o(XDT[8]), .i(CONV_DONE));
buft N91P_13_8 (.i(CREGSEL), .o(XDT[7]), .t(XREG_OUTCS_RD_n));
buft N91P_13_7 (.t(XREG_OUTCS_RD_n), .o(XDT[6]), .i(FECSEL));
buft N91P_13_6 (.t(XREG_OUTCS_RD_n), .o(XDT[5]), .i(LATCH4));
buft N91P_13_5 (.t(XREG_OUTCS_RD_n), .o(XDT[4]), .i(LATCH3));
buft N91P_13_4 (.t(XREG_OUTCS_RD_n), .o(XDT[3]), .i(LATCH2));
buft N91P_13_3 (.t(XREG_OUTCS_RD_n), .o(XDT[2]), .i(LATCH1));
buft N91P_13_2 (.t(XREG_OUTCS_RD_n), .o(XDT[1]), .i(RD_STROBE));
buft N91P_13_1 (.t(XREG_OUTCS_RD_n), .o(XDT[0]), .i(FECBUSY));
buft N88P_13_7 (.i(TAG[4]), .o(XDT[6]), .t(XREG_INCS_RD_n));
buft N88P_13_6 (.t(XREG_INCS_RD_n), .o(XDT[5]), .i(TAG[3]));
buft N88P_13_5 (.t(XREG_INCS_RD_n), .o(XDT[4]), .i(TAG[2]));
buft N88P_13_4 (.t(XREG_INCS_RD_n), .o(XDT[3]), .i(TAG[1]));
buft N88P_13_3 (.t(XREG_INCS_RD_n), .o(XDT[2]), .i(TAG[0]));
buft N88P_13_2 (.t(XREG_INCS_RD_n), .o(XDT[1]), .i(MEMACK2_n));
buft N88P_13_1 (.t(XREG_INCS_RD_n), .o(XDT[0]), .i(CREG_REQ));
buft N111P_13_32 (.i(DAVAIL[32]), .o(XDT[31]), .t(XREG_DAV_RD_n));
buft N111P_13_31 (.t(XREG_DAV_RD_n), .o(XDT[30]), .i(DAVAIL[31]));
buft N111P_13_30 (.t(XREG_DAV_RD_n), .o(XDT[29]), .i(DAVAIL[30]));
buft N111P_13_29 (.t(XREG_DAV_RD_n), .o(XDT[28]), .i(DAVAIL[29]));
buft N111P_13_28 (.t(XREG_DAV_RD_n), .o(XDT[27]), .i(DAVAIL[28]));
buft N111P_13_27 (.t(XREG_DAV_RD_n), .o(XDT[26]), .i(DAVAIL[27]));
buft N111P_13_26 (.t(XREG_DAV_RD_n), .o(XDT[25]), .i(DAVAIL[26]));
buft N111P_13_25 (.t(XREG_DAV_RD_n), .o(XDT[24]), .i(DAVAIL[25]));
buft N111P_13_24 (.t(XREG_DAV_RD_n), .o(XDT[23]), .i(DAVAIL[24]));
buft N111P_13_23 (.t(XREG_DAV_RD_n), .o(XDT[22]), .i(DAVAIL[23]));
buft N111P_13_22 (.t(XREG_DAV_RD_n), .o(XDT[21]), .i(DAVAIL[22]));
buft N111P_13_21 (.t(XREG_DAV_RD_n), .o(XDT[20]), .i(DAVAIL[21]));
buft N111P_13_20 (.t(XREG_DAV_RD_n), .o(XDT[19]), .i(DAVAIL[20]));
buft N111P_13_19 (.t(XREG_DAV_RD_n), .o(XDT[18]), .i(DAVAIL[19]));
buft N111P_13_18 (.t(XREG_DAV_RD_n), .o(XDT[17]), .i(DAVAIL[18]));
buft N111P_13_17 (.t(XREG_DAV_RD_n), .o(XDT[16]), .i(DAVAIL[17]));
buft N111P_13_16 (.t(XREG_DAV_RD_n), .o(XDT[15]), .i(DAVAIL[16]));
buft N111P_13_15 (.t(XREG_DAV_RD_n), .o(XDT[14]), .i(DAVAIL[15]));
buft N111P_13_14 (.t(XREG_DAV_RD_n), .o(XDT[13]), .i(DAVAIL[14]));
buft N111P_13_13 (.t(XREG_DAV_RD_n), .o(XDT[12]), .i(DAVAIL[13]));
buft N111P_13_12 (.t(XREG_DAV_RD_n), .o(XDT[11]), .i(DAVAIL[12]));
buft N111P_13_11 (.t(XREG_DAV_RD_n), .o(XDT[10]), .i(DAVAIL[11]));
buft N111P_13_10 (.t(XREG_DAV_RD_n), .o(XDT[9]), .i(DAVAIL[10]));
buft N111P_13_9 (.t(XREG_DAV_RD_n), .o(XDT[8]), .i(DAVAIL[9]));
buft N111P_13_8 (.t(XREG_DAV_RD_n), .o(XDT[7]), .i(DAVAIL[8]));
buft N111P_13_7 (.t(XREG_DAV_RD_n), .o(XDT[6]), .i(DAVAIL[7]));
buft N111P_13_6 (.t(XREG_DAV_RD_n), .o(XDT[5]), .i(DAVAIL[6]));
buft N111P_13_5 (.t(XREG_DAV_RD_n), .o(XDT[4]), .i(DAVAIL[5]));
buft N111P_13_4 (.t(XREG_DAV_RD_n), .o(XDT[3]), .i(DAVAIL[4]));
buft N111P_13_3 (.t(XREG_DAV_RD_n), .o(XDT[2]), .i(DAVAIL[3]));
buft N111P_13_2 (.t(XREG_DAV_RD_n), .o(XDT[1]), .i(DAVAIL[2]));
buft N111P_13_1 (.t(XREG_DAV_RD_n), .o(XDT[0]), .i(DAVAIL[1]));
aclk N110P_13 (.i(UN_13_ACLK_110P_I), .o(XREG_CDIS_WR));
obuft N4P_6_32 (.i(XDT[31]), .o(BXDT[31]), .t(XREG_RD_n));
obuft N4P_6_31 (.t(XREG_RD_n), .o(BXDT[30]), .i(XDT[30]));
obuft N4P_6_30 (.t(XREG_RD_n), .o(BXDT[29]), .i(XDT[29]));
obuft N4P_6_29 (.t(XREG_RD_n), .o(BXDT[28]), .i(XDT[28]));
obuft N4P_6_28 (.t(XREG_RD_n), .o(BXDT[27]), .i(XDT[27]));
obuft N4P_6_27 (.t(XREG_RD_n), .o(BXDT[26]), .i(XDT[26]));
obuft N4P_6_26 (.t(XREG_RD_n), .o(BXDT[25]), .i(XDT[25]));
obuft N4P_6_25 (.t(XREG_RD_n), .o(BXDT[24]), .i(XDT[24]));
obuft N4P_6_24 (.t(XREG_RD_n), .o(BXDT[23]), .i(XDT[23]));
obuft N4P_6_23 (.t(XREG_RD_n), .o(BXDT[22]), .i(XDT[22]));
obuft N4P_6_22 (.t(XREG_RD_n), .o(BXDT[21]), .i(XDT[21]));
obuft N4P_6_21 (.t(XREG_RD_n), .o(BXDT[20]), .i(XDT[20]));
obuft N4P_6_20 (.t(XREG_RD_n), .o(BXDT[19]), .i(XDT[19]));
obuft N4P_6_19 (.t(XREG_RD_n), .o(BXDT[18]), .i(XDT[18]));
obuft N4P_6_18 (.t(XREG_RD_n), .o(BXDT[17]), .i(XDT[17]));
obuft N4P_6_17 (.t(XREG_RD_n), .o(BXDT[16]), .i(XDT[16]));
obuft N4P_6_16 (.t(XREG_RD_n), .o(BXDT[15]), .i(XDT[15]));
obuft N4P_6_15 (.t(XREG_RD_n), .o(BXDT[14]), .i(XDT[14]));
obuft N4P_6_14 (.t(XREG_RD_n), .o(BXDT[13]), .i(XDT[13]));
obuft N4P_6_13 (.t(XREG_RD_n), .o(BXDT[12]), .i(XDT[12]));
obuft N4P_6_12 (.t(XREG_RD_n), .o(BXDT[11]), .i(XDT[11]));
obuft N4P_6_11 (.t(XREG_RD_n), .o(BXDT[10]), .i(XDT[10]));
obuft N4P_6_10 (.t(XREG_RD_n), .o(BXDT[9]), .i(XDT[9]));
obuft N4P_6_9 (.t(XREG_RD_n), .o(BXDT[8]), .i(XDT[8]));
obuft N4P_6_8 (.t(XREG_RD_n), .o(BXDT[7]), .i(XDT[7]));
obuft N4P_6_7 (.t(XREG_RD_n), .o(BXDT[6]), .i(XDT[6]));
obuft N4P_6_6 (.t(XREG_RD_n), .o(BXDT[5]), .i(XDT[5]));
obuft N4P_6_5 (.t(XREG_RD_n), .o(BXDT[4]), .i(XDT[4]));
obuft N4P_6_4 (.t(XREG_RD_n), .o(BXDT[3]), .i(XDT[3]));
obuft N4P_6_3 (.t(XREG_RD_n), .o(BXDT[2]), .i(XDT[2]));
obuft N4P_6_2 (.t(XREG_RD_n), .o(BXDT[1]), .i(XDT[1]));
obuft N4P_6_1 (.t(XREG_RD_n), .o(BXDT[0]), .i(XDT[0]));
nand4 N137P_5 (.i3(UN_5_NAND4_137P_I3), .o(TAG[2]), .i1(UN_5_NAND4_137P_I1), .i0(UN_5_NAND4_137P_I0), .i2(UN_5_NAND4_137P_I2));
nand4 N136P_5 (.i3(UN_5_NAND4_136P_I3), .o(TAG[1]), .i1(UN_5_NAND4_136P_I1), .i0(UN_5_NAND4_136P_I0), .i2(UN_5_NAND4_136P_I2));
nand4 N135P_5 (.i3(UN_5_NAND4_135P_I3), .o(TAG[0]), .i1(UN_5_NAND4_135P_I1), .i0(UN_5_NAND4_135P_I0), .i2(UN_5_NAND4_135P_I2));
or4 N134P_5 (.i3(EO[3]), .o(DAVAILS), .i1(EO[1]), .i0(EO[0]), .i2(EO[2]));
nor3 N214P_2 (.o(MEMREQ2_n), .i1(REQ2_W2), .i0(REQ2_W1), .i2(REQ2_W3));
and3 N209P_2 (.o(REQ2_W2), .i1(MEMACK2_n), .i0(CAD_EN_n), .i2(UN_2_AND3_209P_I2));
and3 N208P_2 (.o(REQ2_W1), .i1(UN_2_AND3_208P_I1), .i0(MEMACK2_n), .i2(UN_2_AND3_208P_I2));
ofd N150P_5_5 (.q(BTAG[4]), .d(TAG[4]), .c(CHIP_SEL_EN), .gr(RESET_n));
ofd N150P_5_4 (.c(CHIP_SEL_EN), .d(TAG[3]), .q(BTAG[3]), .gr(RESET_n));
ofd N150P_5_3 (.c(CHIP_SEL_EN), .d(TAG[2]), .q(BTAG[2]), .gr(RESET_n));
ofd N150P_5_2 (.c(CHIP_SEL_EN), .d(TAG[1]), .q(BTAG[1]), .gr(RESET_n));
ofd N150P_5_1 (.c(CHIP_SEL_EN), .d(TAG[0]), .q(BTAG[0]), .gr(RESET_n));
obuf N230P_1_4 (.i(LATCH4), .o(BLATCH[4]));
obuf N230P_1_3 (.o(BLATCH[3]), .i(LATCH3));
obuf N230P_1_2 (.o(BLATCH[2]), .i(LATCH2));
obuf N230P_1_1 (.o(BLATCH[1]), .i(LATCH1));
obuf N2P_10 (.i(DOUT), .o(SDOUT));
obuf N3P_10 (.i(SM2), .o(M2));
obuf N168P_3 (.i(CONV_DONE), .o(BCONV_DONE));
obuf N156P_3 (.i(ADC_CONVERT_n), .o(BADC_CONVERT_n));
obuf N195P_2 (.i(MEMREQ2_n), .o(BMEMREQ2_n));
obuf N265P_1 (.i(CREGSEL), .o(BCREGSEL));
obuf N245P_1 (.i(RD_STROBE), .o(BRD_STROBE));
obuf N242P_1 (.i(CHOLD_n), .o(BCHOLD_n));
obuf N236P_1 (.i(CAD_EN), .o(BCAD_EN));
obuf N234P_1 (.i(CHIP_SEL_EN), .o(BCHIP_SEL_EN));
obuf N228P_1 (.i(FECBUSY), .o(BFECBUSY));
obuf N212P_2_3 (.i(ENW1_n), .o(BN_ENW[3]));
obuf N212P_2_2 (.o(BN_ENW[2]), .i(ENW2_n));
obuf N212P_2_1 (.o(BN_ENW[1]), .i(ENW3_n));
ibuf N3P_6_32 (.i(BDAVAIL[32]), .o(DAVAIL[32]));
ibuf N3P_6_31 (.o(DAVAIL[31]), .i(BDAVAIL[31]));
ibuf N3P_6_30 (.o(DAVAIL[30]), .i(BDAVAIL[30]));
ibuf N3P_6_29 (.o(DAVAIL[29]), .i(BDAVAIL[29]));
ibuf N3P_6_28 (.o(DAVAIL[28]), .i(BDAVAIL[28]));
ibuf N3P_6_27 (.o(DAVAIL[27]), .i(BDAVAIL[27]));
ibuf N3P_6_26 (.o(DAVAIL[26]), .i(BDAVAIL[26]));
ibuf N3P_6_25 (.o(DAVAIL[25]), .i(BDAVAIL[25]));
ibuf N3P_6_24 (.o(DAVAIL[24]), .i(BDAVAIL[24]));
ibuf N3P_6_23 (.o(DAVAIL[23]), .i(BDAVAIL[23]));
ibuf N3P_6_22 (.o(DAVAIL[22]), .i(BDAVAIL[22]));
ibuf N3P_6_21 (.o(DAVAIL[21]), .i(BDAVAIL[21]));
ibuf N3P_6_20 (.o(DAVAIL[20]), .i(BDAVAIL[20]));
ibuf N3P_6_19 (.o(DAVAIL[19]), .i(BDAVAIL[19]));
ibuf N3P_6_18 (.o(DAVAIL[18]), .i(BDAVAIL[18]));
ibuf N3P_6_17 (.o(DAVAIL[17]), .i(BDAVAIL[17]));
ibuf N3P_6_16 (.o(DAVAIL[16]), .i(BDAVAIL[16]));
ibuf N3P_6_15 (.o(DAVAIL[15]), .i(BDAVAIL[15]));
ibuf N3P_6_14 (.o(DAVAIL[14]), .i(BDAVAIL[14]));
ibuf N3P_6_13 (.o(DAVAIL[13]), .i(BDAVAIL[13]));
ibuf N3P_6_12 (.o(DAVAIL[12]), .i(BDAVAIL[12]));
ibuf N3P_6_11 (.o(DAVAIL[11]), .i(BDAVAIL[11]));
ibuf N3P_6_10 (.o(DAVAIL[10]), .i(BDAVAIL[10]));
ibuf N3P_6_9 (.o(DAVAIL[9]), .i(BDAVAIL[9]));
ibuf N3P_6_8 (.o(DAVAIL[8]), .i(BDAVAIL[8]));
ibuf N3P_6_7 (.o(DAVAIL[7]), .i(BDAVAIL[7]));
ibuf N3P_6_6 (.o(DAVAIL[6]), .i(BDAVAIL[6]));
ibuf N3P_6_5 (.o(DAVAIL[5]), .i(BDAVAIL[5]));
ibuf N3P_6_4 (.o(DAVAIL[4]), .i(BDAVAIL[4]));
ibuf N3P_6_3 (.o(DAVAIL[3]), .i(BDAVAIL[3]));
ibuf N3P_6_2 (.o(DAVAIL[2]), .i(BDAVAIL[2]));
ibuf N3P_6_1 (.o(DAVAIL[1]), .i(BDAVAIL[1]));
ibuf N6P_6_32 (.i(BXDT[31]), .o(XD[31]));
ibuf N6P_6_31 (.o(XD[30]), .i(BXDT[30]));
ibuf N6P_6_30 (.o(XD[29]), .i(BXDT[29]));
ibuf N6P_6_29 (.o(XD[28]), .i(BXDT[28]));
ibuf N6P_6_28 (.o(XD[27]), .i(BXDT[27]));
ibuf N6P_6_27 (.o(XD[26]), .i(BXDT[26]));
ibuf N6P_6_26 (.o(XD[25]), .i(BXDT[25]));
ibuf N6P_6_25 (.o(XD[24]), .i(BXDT[24]));
ibuf N6P_6_24 (.o(XD[23]), .i(BXDT[23]));
ibuf N6P_6_23 (.o(XD[22]), .i(BXDT[22]));
ibuf N6P_6_22 (.o(XD[21]), .i(BXDT[21]));
ibuf N6P_6_21 (.o(XD[20]), .i(BXDT[20]));
ibuf N6P_6_20 (.o(XD[19]), .i(BXDT[19]));
ibuf N6P_6_19 (.o(XD[18]), .i(BXDT[18]));
ibuf N6P_6_18 (.o(XD[17]), .i(BXDT[17]));
ibuf N6P_6_17 (.o(XD[16]), .i(BXDT[16]));
ibuf N6P_6_16 (.o(XD[15]), .i(BXDT[15]));
ibuf N6P_6_15 (.o(XD[14]), .i(BXDT[14]));
ibuf N6P_6_14 (.o(XD[13]), .i(BXDT[13]));
ibuf N6P_6_13 (.o(XD[12]), .i(BXDT[12]));
ibuf N6P_6_12 (.o(XD[11]), .i(BXDT[11]));
ibuf N6P_6_11 (.o(XD[10]), .i(BXDT[10]));
ibuf N6P_6_10 (.o(XD[9]), .i(BXDT[9]));
ibuf N6P_6_9 (.o(XD[8]), .i(BXDT[8]));
ibuf N6P_6_8 (.o(XD[7]), .i(BXDT[7]));
ibuf N6P_6_7 (.o(XD[6]), .i(BXDT[6]));
ibuf N6P_6_6 (.o(XD[5]), .i(BXDT[5]));
ibuf N6P_6_5 (.o(XD[4]), .i(BXDT[4]));
ibuf N6P_6_4 (.o(XD[3]), .i(BXDT[3]));
ibuf N6P_6_3 (.o(XD[2]), .i(BXDT[2]));
ibuf N6P_6_2 (.o(XD[1]), .i(BXDT[1]));
ibuf N6P_6_1 (.o(XD[0]), .i(BXDT[0]));
ibuf N26P_13 (.i(BXREG_WR_n), .o(XREG_WR_n));
ibuf N27P_13 (.i(BXREG_RD_n), .o(XREG_RD_n));
ibuf N6P_10 (.i(SDIN), .o(DIN));
ibuf N185P_2 (.i(BMEMACK2_n), .o(MEMACK2_n));
ibuf N257P_1 (.i(BCLKA), .o(CLKA));
ibuf N221P_1 (.i(BSEQ_RESET), .o(SEQ_RESET));
ibuf N220P_1 (.i(BCREG_REQ), .o(CREG_REQ));
ibuf N35P_13_3 (.i(BXREG_SEL[2]), .o(XREG_SEL[2]));
ibuf N35P_13_2 (.o(XREG_SEL[1]), .i(BXREG_SEL[1]));
ibuf N35P_13_1 (.o(XREG_SEL[0]), .i(BXREG_SEL[0]));
gclk N218P_1 (.i(BCLK), .o(CLK));
nand2 N7P_6_32 (.o(DAVM_[32]), .i1(DAVAIL[32]), .i0(CHIP_MASK[32]));
nand2 N7P_6_31 (.i0(CHIP_MASK[31]), .i1(DAVAIL[31]), .o(DAVM_[31]));
nand2 N7P_6_30 (.i0(CHIP_MASK[30]), .i1(DAVAIL[30]), .o(DAVM_[30]));
nand2 N7P_6_29 (.i0(CHIP_MASK[29]), .i1(DAVAIL[29]), .o(DAVM_[29]));
nand2 N7P_6_28 (.i0(CHIP_MASK[28]), .i1(DAVAIL[28]), .o(DAVM_[28]));
nand2 N7P_6_27 (.i0(CHIP_MASK[27]), .i1(DAVAIL[27]), .o(DAVM_[27]));
nand2 N7P_6_26 (.i0(CHIP_MASK[26]), .i1(DAVAIL[26]), .o(DAVM_[26]));
nand2 N7P_6_25 (.i0(CHIP_MASK[25]), .i1(DAVAIL[25]), .o(DAVM_[25]));
nand2 N7P_6_24 (.i0(CHIP_MASK[24]), .i1(DAVAIL[24]), .o(DAVM_[24]));
nand2 N7P_6_23 (.i0(CHIP_MASK[23]), .i1(DAVAIL[23]), .o(DAVM_[23]));
nand2 N7P_6_22 (.i0(CHIP_MASK[22]), .i1(DAVAIL[22]), .o(DAVM_[22]));
nand2 N7P_6_21 (.i0(CHIP_MASK[21]), .i1(DAVAIL[21]), .o(DAVM_[21]));
nand2 N7P_6_20 (.i0(CHIP_MASK[20]), .i1(DAVAIL[20]), .o(DAVM_[20]));
nand2 N7P_6_19 (.i0(CHIP_MASK[19]), .i1(DAVAIL[19]), .o(DAVM_[19]));
nand2 N7P_6_18 (.i0(CHIP_MASK[18]), .i1(DAVAIL[18]), .o(DAVM_[18]));
nand2 N7P_6_17 (.i0(CHIP_MASK[17]), .i1(DAVAIL[17]), .o(DAVM_[17]));
nand2 N7P_6_16 (.i0(CHIP_MASK[16]), .i1(DAVAIL[16]), .o(DAVM_[16]));
nand2 N7P_6_15 (.i0(CHIP_MASK[15]), .i1(DAVAIL[15]), .o(DAVM_[15]));
nand2 N7P_6_14 (.i0(CHIP_MASK[14]), .i1(DAVAIL[14]), .o(DAVM_[14]));
nand2 N7P_6_13 (.i0(CHIP_MASK[13]), .i1(DAVAIL[13]), .o(DAVM_[13]));
nand2 N7P_6_12 (.i0(CHIP_MASK[12]), .i1(DAVAIL[12]), .o(DAVM_[12]));
nand2 N7P_6_11 (.i0(CHIP_MASK[11]), .i1(DAVAIL[11]), .o(DAVM_[11]));
nand2 N7P_6_10 (.i0(CHIP_MASK[10]), .i1(DAVAIL[10]), .o(DAVM_[10]));
nand2 N7P_6_9 (.i0(CHIP_MASK[9]), .i1(DAVAIL[9]), .o(DAVM_[9]));
nand2 N7P_6_8 (.i0(CHIP_MASK[8]), .i1(DAVAIL[8]), .o(DAVM_[8]));
nand2 N7P_6_7 (.i0(CHIP_MASK[7]), .i1(DAVAIL[7]), .o(DAVM_[7]));
nand2 N7P_6_6 (.i0(CHIP_MASK[6]), .i1(DAVAIL[6]), .o(DAVM_[6]));
nand2 N7P_6_5 (.i0(CHIP_MASK[5]), .i1(DAVAIL[5]), .o(DAVM_[5]));
nand2 N7P_6_4 (.i0(CHIP_MASK[4]), .i1(DAVAIL[4]), .o(DAVM_[4]));
nand2 N7P_6_3 (.i0(CHIP_MASK[3]), .i1(DAVAIL[3]), .o(DAVM_[3]));
nand2 N7P_6_2 (.i0(CHIP_MASK[2]), .i1(DAVAIL[2]), .o(DAVM_[2]));
nand2 N7P_6_1 (.i0(CHIP_MASK[1]), .i1(DAVAIL[1]), .o(DAVM_[1]));
nand2 N181P_2 (.o(MEMCLR_n), .i1(WRITEDONE_n), .i0(SEQ_RESET_n));
nand2 N167P_2 (.o(ENW2_n), .i1(REQ2_W2), .i0(ENW3_n));
nand2 N208P_1 (.o(UN_1_FDC_183P_CLR), .i1(UN_1_NAND2_208P_I1), .i0(SEQ_RESET));
nand2 N206P_1 (.i0(XVDD), .o(UN_1_FDC_205P_CLR), .i1(CDONE_n));
nor2 N1P_6_32 (.o(CHIP_MASK[32]), .i1(LAST_SELECTED_[32]), .i0(CDIS[32]));
nor2 N1P_6_31 (.i0(CDIS[31]), .i1(LAST_SELECTED_[31]), .o(CHIP_MASK[31]));
nor2 N1P_6_30 (.i0(CDIS[30]), .i1(LAST_SELECTED_[30]), .o(CHIP_MASK[30]));
nor2 N1P_6_29 (.i0(CDIS[29]), .i1(LAST_SELECTED_[29]), .o(CHIP_MASK[29]));
nor2 N1P_6_28 (.i0(CDIS[28]), .i1(LAST_SELECTED_[28]), .o(CHIP_MASK[28]));
nor2 N1P_6_27 (.i0(CDIS[27]), .i1(LAST_SELECTED_[27]), .o(CHIP_MASK[27]));
nor2 N1P_6_26 (.i0(CDIS[26]), .i1(LAST_SELECTED_[26]), .o(CHIP_MASK[26]));
nor2 N1P_6_25 (.i0(CDIS[25]), .i1(LAST_SELECTED_[25]), .o(CHIP_MASK[25]));
nor2 N1P_6_24 (.i0(CDIS[24]), .i1(LAST_SELECTED_[24]), .o(CHIP_MASK[24]));
nor2 N1P_6_23 (.i0(CDIS[23]), .i1(LAST_SELECTED_[23]), .o(CHIP_MASK[23]));
nor2 N1P_6_22 (.i0(CDIS[22]), .i1(LAST_SELECTED_[22]), .o(CHIP_MASK[22]));
nor2 N1P_6_21 (.i0(CDIS[21]), .i1(LAST_SELECTED_[21]), .o(CHIP_MASK[21]));
nor2 N1P_6_20 (.i0(CDIS[20]), .i1(LAST_SELECTED_[20]), .o(CHIP_MASK[20]));
nor2 N1P_6_19 (.i0(CDIS[19]), .i1(LAST_SELECTED_[19]), .o(CHIP_MASK[19]));
nor2 N1P_6_18 (.i0(CDIS[18]), .i1(LAST_SELECTED_[18]), .o(CHIP_MASK[18]));
nor2 N1P_6_17 (.i0(CDIS[17]), .i1(LAST_SELECTED_[17]), .o(CHIP_MASK[17]));
nor2 N1P_6_16 (.i0(CDIS[16]), .i1(LAST_SELECTED_[16]), .o(CHIP_MASK[16]));
nor2 N1P_6_15 (.i0(CDIS[15]), .i1(LAST_SELECTED_[15]), .o(CHIP_MASK[15]));
nor2 N1P_6_14 (.i0(CDIS[14]), .i1(LAST_SELECTED_[14]), .o(CHIP_MASK[14]));
nor2 N1P_6_13 (.i0(CDIS[13]), .i1(LAST_SELECTED_[13]), .o(CHIP_MASK[13]));
nor2 N1P_6_12 (.i0(CDIS[12]), .i1(LAST_SELECTED_[12]), .o(CHIP_MASK[12]));
nor2 N1P_6_11 (.i0(CDIS[11]), .i1(LAST_SELECTED_[11]), .o(CHIP_MASK[11]));
nor2 N1P_6_10 (.i0(CDIS[10]), .i1(LAST_SELECTED_[10]), .o(CHIP_MASK[10]));
nor2 N1P_6_9 (.i0(CDIS[9]), .i1(LAST_SELECTED_[9]), .o(CHIP_MASK[9]));
nor2 N1P_6_8 (.i0(CDIS[8]), .i1(LAST_SELECTED_[8]), .o(CHIP_MASK[8]));
nor2 N1P_6_7 (.i0(CDIS[7]), .i1(LAST_SELECTED_[7]), .o(CHIP_MASK[7]));
nor2 N1P_6_6 (.i0(CDIS[6]), .i1(LAST_SELECTED_[6]), .o(CHIP_MASK[6]));
nor2 N1P_6_5 (.i0(CDIS[5]), .i1(LAST_SELECTED_[5]), .o(CHIP_MASK[5]));
nor2 N1P_6_4 (.i0(CDIS[4]), .i1(LAST_SELECTED_[4]), .o(CHIP_MASK[4]));
nor2 N1P_6_3 (.i0(CDIS[3]), .i1(LAST_SELECTED_[3]), .o(CHIP_MASK[3]));
nor2 N1P_6_2 (.i0(CDIS[2]), .i1(LAST_SELECTED_[2]), .o(CHIP_MASK[2]));
nor2 N1P_6_1 (.i0(CDIS[1]), .i1(LAST_SELECTED_[1]), .o(CHIP_MASK[1]));
nor2 N193P_1 (.o(UN_1_FDC_191P_D), .i1(FECSTART), .i0(CHOLD_n));
inv N149P_5 (.i(UN_5_INV_149P_I), .o(TAG[3]));
inv N148P_5 (.i(UN_5_INV_148P_I), .o(TAG[4]));
inv N133P_5 (.i(DAVAILS), .o(DAVAILS_n));
inv N77P_4 (.i(TAG[4]), .o(UN_4_INV_77P_O));
inv N76P_4 (.i(TAG[3]), .o(UN_4_INV_76P_O));
inv N175P_3 (.i(UN_3_FDC_133P_Q), .o(UN_3_FDC_133P_D));
inv N174P_3 (.i(UN_3_FDC_128P_Q), .o(UN_3_FDC_136P_C));
inv N172P_3 (.i(UN_3_FDC_139P_Q), .o(UN_3_FDC_128P_C));
inv N171P_3 (.i(UN_3_FDC_144P_Q), .o(UN_3_FDC_142P_C));
inv N173P_3 (.i(UN_3_FDC_142P_Q), .o(UN_3_FDC_142P_D));
inv N162P_3 (.i(UN_3_FDC_166P_Q), .o(CAD_EN_START_n));
inv N157P_3 (.i(UN_3_FDC_127P_Q), .o(UN_3_FDC_126P_D));
inv N135P_3 (.i(UN_3_FDC_136P_Q), .o(UN_3_FDC_133P_C));
inv N125P_3 (.i(ADC_CONVERT), .o(ADC_CONVERT_n));
inv N175P_2 (.i(UN_2_AND3_208P_I1), .o(MEMWR2_n));
inv N174P_2 (.i(MEMACK2_n), .o(UN_2_FDC_171P_C));
inv N170P_2 (.i(UN_2_AND3_209P_I2), .o(UN_2_AND3_208P_I2));
inv N169P_2 (.i(UN_2_FDC_171P_Q), .o(WRITEDONE_n));
inv N166P_2 (.i(REQ2_W1), .o(ENW1_n));
inv N165P_2 (.i(REQ2_W3), .o(ENW3_n));
inv N164P_2 (.i(SEQ_RESET), .o(SEQ_RESET_n));
inv N196P_2 (.i(CAD_EN), .o(CAD_EN_n));
inv N261P_1 (.i(CDONE), .o(CDONE_n));
inv N260P_1 (.i(UN_1_FDC_205P_Q), .o(CHOLD_n));
inv N258P_1 (.i(CLKA), .o(CLKA_n));
inv N212P_1 (.i(UN_1_FDC_213P_Q), .o(UN_1_INV_212P_O));
inv N210P_1 (.i(CREGSEL_n), .o(CREGSEL));
inv N209P_1 (.i(FECSEL_n), .o(FECSEL));
inv N194P_1 (.i(CLK), .o(CLK_n));
inv N185P_1 (.i(FECSEL_n), .o(CREGSEL_n));
inv N184P_1 (.i(UN_1_FDC_183P_Q), .o(UN_1_INV_184P_O));
and2 N210P_2 (.o(REQ2_W3), .i1(UN_2_AND2_210P_I1), .i0(MEMACK2_n));
and2 N263P_1 (.o(UN_1_AND2_263P_O), .i1(UN_1_AND2_182P_O), .i0(CHOLD_n));
and2 N262P_1 (.o(UN_1_AND2_262P_O), .i1(RD_STROBE), .i0(LATCH4));
and2 N187P_1 (.o(UN_1_AND2_187P_O), .i1(DAVAILS), .i0(CREGSEL_n));
and2 N182P_1 (.o(UN_1_AND2_182P_O), .i1(DAVAILS), .i0(MEMWR2_n));
or2 N132P_5 (.o(DAV_n), .i1(DAVAILS_n), .i0(SEQ_RESET));
or2 N153P_3 (.o(UN_3_FDC_132P_CLR), .i1(UN_3_FDC_131P_Q), .i0(SEQ_RESET));
or2 N145P_3 (.o(UN_3_FDC_142P_CLR), .i1(SEQ_RESET), .i0(CAD_EN_START_n));
or2 N141P_3 (.o(CONV_DONE), .i1(UN_3_FDC_131P_D), .i0(SEQ_RESET));
or2 N176P_2 (.o(UN_2_FDC_180P_D), .i1(UN_2_AND3_208P_I1), .i0(CREGSEL_n));
or2 N215P_1 (.o(RD_STROBE), .i1(CLKA_n), .i0(UN_1_INV_212P_O));
or2 N196P_1 (.o(UN_1_FDC_192P_D), .i1(FECSTART), .i0(UN_1_AND2_263P_O));
or2 N195P_1 (.o(UPSTART), .i1(FECSTART), .i0(FECSEL_n));
or2 N190P_1 (.o(UN_1_FDC_183P_D), .i1(UN_1_FDC_183P_Q), .i0(FECSTART));
or2 N189P_1 (.o(FECBUSY), .i1(UN_1_AND2_187P_O), .i0(UN_1_FDC_183P_Q));
or2 N188P_1 (.o(UN_1_NAND2_208P_I1), .i1(UN_1_INV_184P_O), .i0(WRITEDONE_n));
or2 N180P_1 (.o(CDONE), .i1(CONV_DONE), .i0(SEQ_RESET));
endmodule
`uselib

module sequencer32_globals();

wire GR;
endmodule

