/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from seq96newt.xcd on Fri Jul  5 16:05:42 1996 */
/* PART 3064APQ160-6 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module seq96newt
(SQXREG_WR_n, SQXREG_SEL, SQXREG_RD_n, SQTAG, SQRD_STROBE_n, SQMEMORY_REQUEST_n, SQMEMORY_ACK_n, SQLATCH, SQFECBUSY, SQENW_, SQDAV32OR, SQDAV, SQD, SQCREG_SEL, SQCREG_REQ, SQCONVERT_START_n, SQCLK, SQCHOLD_n, SQCHIP_SEL_EN, SQCADD_ENABLE, SQADC_BUSY_n, SPAREOUT, SPAREIN, SDOUT, SDIN, M2, RESET_n, ADC_DONE, RDATA_n, RTRIG, PROGRAM_n, CCLK, PWRDWN_n);
   input SQXREG_WR_n;
   input [2:0] SQXREG_SEL;
   input SQXREG_RD_n;
   output [4:0] SQTAG;
   output SQRD_STROBE_n;
   output SQMEMORY_REQUEST_n;
   input SQMEMORY_ACK_n;
   output [4:1] SQLATCH;
   output SQFECBUSY;
   output [3:1] SQENW_;
   output SQDAV32OR;
   input [32:1] SQDAV;
   inout [31:0] SQD;
   output SQCREG_SEL;
   input SQCREG_REQ;
   output SQCONVERT_START_n;
   input SQCLK;
   output SQCHOLD_n;
   output SQCHIP_SEL_EN;
   output SQCADD_ENABLE;
   input SQADC_BUSY_n;
   output [2:0] SPAREOUT;
   input [2:0] SPAREIN;
   output SDOUT;
   input SDIN;
   output M2;
   input RESET_n;
   output ADC_DONE;
   output RDATA_n;
   input RTRIG;
   input PROGRAM_n;
   input CCLK;
   input PWRDWN_n;
wire [31:0] N47P_1_DOUT;
wire [31:0] N47P_1_DIN;
wire [0:0] N31P_1_4P_1_19P_1_I18_1_I7_1_QD;
wire [0:0] N31P_1_4P_1_19P_1_I18_1_I7_1_A1;
wire [0:0] N31P_1_4P_1_19P_1_I18_1_D_S;
wire [0:0] N31P_1_4P_1_19P_1_I15_1_I7_1_QD;
wire [0:0] N31P_1_4P_1_19P_1_I15_1_I7_1_A1;
wire [0:0] N31P_1_4P_1_19P_1_I15_1_D_S;
wire [0:0] N31P_1_4P_1_19P_1_I14_1_I7_1_QD;
wire [0:0] N31P_1_4P_1_19P_1_I14_1_I7_1_A1;
wire [0:0] N31P_1_4P_1_19P_1_I14_1_D_S;
wire [0:0] N31P_1_4P_1_19P_1_I13_1_I7_1_QD;
wire [0:0] N31P_1_4P_1_19P_1_I13_1_I7_1_A1;
wire [0:0] N31P_1_4P_1_19P_1_I13_1_D_S;
wire [3:1] N31P_1_4P_1_STAGE;
wire [3:0] N31P_1_4P_1_S;
wire [3:0] N31P_1_4P_1_C;
wire [0:0] N31P_1_2P_1_83P_1_I34_1_TQ;
wire [0:0] N31P_1_2P_1_83P_1_I30_1_TQ;
wire [0:0] N31P_1_2P_1_83P_1_I28_1_TQ;
wire [0:0] N31P_1_2P_1_83P_1_I26_1_TQ;
wire [0:0] N31P_1_2P_1_83P_1_I23_1_TQ;
wire [0:0] N31P_1_2P_1_83P_1_I20_1_TQ;
wire [0:0] N31P_1_2P_1_83P_1_I18_1_TQ;
wire [0:0] N31P_1_2P_1_83P_1_I15_1_TQ;
wire [5:0] N31P_1_2P_1_WAIT;
wire [4:1] N31P_1_2P_1_STROBE;
wire [7:0] N31P_1_2P_1_STATES;
wire [0:0] N6P_1_17P_1_I34_1_TQ;
wire [0:0] N6P_1_17P_1_I30_1_TQ;
wire [0:0] N6P_1_17P_1_I28_1_TQ;
wire [0:0] N6P_1_17P_1_I26_1_TQ;
wire [0:0] N6P_1_17P_1_I23_1_TQ;
wire [0:0] N6P_1_17P_1_I20_1_TQ;
wire [0:0] N6P_1_17P_1_I18_1_TQ;
wire [0:0] N6P_1_17P_1_I15_1_TQ;
wire [0:0] N6P_1_5P_2_I47;
wire [0:0] N6P_1_4P_2_I47;
wire [0:0] N6P_1_4P_1_I47;
wire [0:0] N6P_1_3P_2_I47;
wire [0:0] N6P_1_3P_1_I47;
wire [0:0] N6P_1_2P_1_I47;
wire [0:0] N6P_1_1P_2_I47;
wire [0:0] N6P_1_1P_1_I47;
wire [32:1] N6P_1_SELECT;
wire [7:0] N6P_1_FULL_TAG;
wire [32:1] N6P_1_CHECK;
wire [2:0] UN_1_AND2_82P_O;
wire [2:0] UN_1_AND2_82P_I0;
wire [4:0] TAG;
wire [2:0] REG_SEL;
wire [4:1] LATCH;
wire [3:1] ENW_;
wire [32:1] DAV;
wire [32:1] CHIP_DISABLE;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/preprod_board/fec32m/develop/seq96newt/verilog_lib/seq96newt.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

fdce N71P_1_I4_1 (.d(GET_DATA), .q(UN_1_FD_1_71P_Q), .c(N71P_1_CB), .ce(XVDD), .clr(XGND), .gr(RESET_n));
inv N71P_1_I5_1 (.i(CLKD2), .o(N71P_1_CB));
or5 N6P_1_1P_2_I10_1 (.i4(N6P_1_1P_2_I47[0]), .i2(DAV[19]), .i3(DAV[20]), .o(N6P_1_UN_2_OR4_2P_I2), .i0(DAV[17]), .i1(DAV[18]));
or4 N6P_1_1P_2_I13_1 (.i2(DAV[23]), .i3(DAV[24]), .o(N6P_1_1P_2_I47[0]), .i0(DAV[21]), .i1(DAV[22]));
or5 N6P_1_5P_2_I10_1 (.i4(N6P_1_5P_2_I47[0]), .i2(DAV[11]), .i3(DAV[12]), .o(N6P_1_UN_2_OR4_2P_I1), .i0(DAV[9]), .i1(DAV[10]));
or4 N6P_1_5P_2_I13_1 (.i2(DAV[15]), .i3(DAV[16]), .o(N6P_1_5P_2_I47[0]), .i0(DAV[13]), .i1(DAV[14]));
or5 N6P_1_4P_2_I10_1 (.i4(N6P_1_4P_2_I47[0]), .i2(DAV[3]), .i3(DAV[4]), .o(N6P_1_UN_2_OR4_2P_I0), .i0(DAV[1]), .i1(DAV[2]));
or4 N6P_1_4P_2_I13_1 (.i2(DAV[7]), .i3(DAV[8]), .o(N6P_1_4P_2_I47[0]), .i0(DAV[5]), .i1(DAV[6]));
or5 N6P_1_3P_2_I10_1 (.i4(N6P_1_3P_2_I47[0]), .i2(DAV[27]), .i3(DAV[28]), .o(N6P_1_UN_2_OR4_2P_I3), .i0(DAV[25]), .i1(DAV[26]));
or4 N6P_1_3P_2_I13_1 (.i2(DAV[31]), .i3(DAV[32]), .o(N6P_1_3P_2_I47[0]), .i0(DAV[29]), .i1(DAV[30]));
or5 N6P_1_1P_1_I10_1 (.i4(N6P_1_1P_1_I47[0]), .i2(N6P_1_SELECT[6]), .i3(N6P_1_SELECT[5]), .o(N6P_1_UN_1_OR4_5P_I3), .i0(N6P_1_SELECT[8]), .i1(N6P_1_SELECT[7]));
or4 N6P_1_1P_1_I13_1 (.i2(N6P_1_SELECT[2]), .i3(N6P_1_SELECT[1]), .o(N6P_1_1P_1_I47[0]), .i0(N6P_1_SELECT[4]), .i1(N6P_1_SELECT[3]));
or5 N6P_1_2P_1_I10_1 (.i4(N6P_1_2P_1_I47[0]), .i2(N6P_1_SELECT[14]), .i3(N6P_1_SELECT[13]), .o(N6P_1_UN_1_OR4_5P_I2), .i0(N6P_1_SELECT[16]), .i1(N6P_1_SELECT[15]));
or4 N6P_1_2P_1_I13_1 (.i2(N6P_1_SELECT[10]), .i3(N6P_1_SELECT[9]), .o(N6P_1_2P_1_I47[0]), .i0(N6P_1_SELECT[12]), .i1(N6P_1_SELECT[11]));
or5 N6P_1_4P_1_I10_1 (.i4(N6P_1_4P_1_I47[0]), .i2(N6P_1_SELECT[30]), .i3(N6P_1_SELECT[29]), .o(N6P_1_UN_1_OR4_5P_I0), .i0(N6P_1_SELECT[32]), .i1(N6P_1_SELECT[31]));
or4 N6P_1_4P_1_I13_1 (.i2(N6P_1_SELECT[26]), .i3(N6P_1_SELECT[25]), .o(N6P_1_4P_1_I47[0]), .i0(N6P_1_SELECT[28]), .i1(N6P_1_SELECT[27]));
or5 N6P_1_3P_1_I10_1 (.i4(N6P_1_3P_1_I47[0]), .i2(N6P_1_SELECT[22]), .i3(N6P_1_SELECT[21]), .o(N6P_1_UN_1_OR4_5P_I1), .i0(N6P_1_SELECT[24]), .i1(N6P_1_SELECT[23]));
or4 N6P_1_3P_1_I13_1 (.i2(N6P_1_SELECT[18]), .i3(N6P_1_SELECT[17]), .o(N6P_1_3P_1_I47[0]), .i0(N6P_1_SELECT[20]), .i1(N6P_1_SELECT[19]));
fdce N6P_1_62P_1_I6_1_5 (.d(N6P_1_FULL_TAG[5]), .q(TAG[4]), .c(DATA_AVAILABLE), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N6P_1_62P_1_I6_1_4 (.clr(XGND), .ce(XVDD), .c(DATA_AVAILABLE), .q(TAG[3]), .d(N6P_1_FULL_TAG[4]), .gr(RESET_n));
fdce N6P_1_62P_1_I6_1_3 (.clr(XGND), .ce(XVDD), .c(DATA_AVAILABLE), .q(TAG[2]), .d(N6P_1_FULL_TAG[3]), .gr(RESET_n));
fdce N6P_1_62P_1_I6_1_2 (.clr(XGND), .ce(XVDD), .c(DATA_AVAILABLE), .q(TAG[1]), .d(N6P_1_FULL_TAG[2]), .gr(RESET_n));
fdce N6P_1_62P_1_I6_1_1 (.clr(XGND), .ce(XVDD), .c(DATA_AVAILABLE), .q(TAG[0]), .d(N6P_1_FULL_TAG[1]), .gr(RESET_n));
and5b4 N6P_1_19P_1_I33_1 (.i4(N6P_1_FULL_TAG[5]), .i3(N6P_1_FULL_TAG[2]), .i2(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[17]), .i1(N6P_1_FULL_TAG[4]), .i0(N6P_1_FULL_TAG[3]));
and5b1 N6P_1_19P_1_I39_1 (.i4(N6P_1_FULL_TAG[5]), .i3(N6P_1_FULL_TAG[2]), .i2(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[24]), .i0(N6P_1_FULL_TAG[4]), .i1(N6P_1_FULL_TAG[3]));
and5b1 N6P_1_19P_1_I30_1 (.i4(N6P_1_FULL_TAG[5]), .i3(N6P_1_FULL_TAG[2]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[28]), .i0(N6P_1_FULL_TAG[3]), .i1(N6P_1_FULL_TAG[1]));
and5b1 N6P_1_19P_1_I29_1 (.i4(N6P_1_FULL_TAG[5]), .i3(N6P_1_FULL_TAG[3]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[30]), .i0(N6P_1_FULL_TAG[2]), .i1(N6P_1_FULL_TAG[1]));
and5b1 N6P_1_19P_1_I25_1 (.i4(N6P_1_FULL_TAG[5]), .i3(N6P_1_FULL_TAG[3]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[31]), .i0(N6P_1_FULL_TAG[1]), .i1(N6P_1_FULL_TAG[2]));
and5b3 N6P_1_19P_1_I37_1 (.i4(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[3]), .i3(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[25]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[2]));
and5b3 N6P_1_19P_1_I35_1 (.i4(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[4]), .i3(N6P_1_FULL_TAG[3]), .o(N6P_1_CHECK[21]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[2]));
and5b3 N6P_1_19P_1_I34_1 (.i4(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[3]), .i3(N6P_1_FULL_TAG[2]), .o(N6P_1_CHECK[19]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[4]));
and5b3 N6P_1_19P_1_I23_1 (.i4(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[4]), .i3(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[18]), .i1(N6P_1_FULL_TAG[2]), .i0(N6P_1_FULL_TAG[3]));
and5b2 N6P_1_19P_1_I36_1 (.i4(N6P_1_FULL_TAG[3]), .i3(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[29]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[2]));
and5b2 N6P_1_19P_1_I31_1 (.i4(N6P_1_FULL_TAG[2]), .i3(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[27]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[3]));
and5b2 N6P_1_19P_1_I32_1 (.i4(N6P_1_FULL_TAG[1]), .i3(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[26]), .i1(N6P_1_FULL_TAG[2]), .i0(N6P_1_FULL_TAG[3]));
and5b2 N6P_1_19P_1_I28_1 (.i4(N6P_1_FULL_TAG[2]), .i3(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[3]), .o(N6P_1_CHECK[23]), .i1(N6P_1_FULL_TAG[4]), .i0(N6P_1_FULL_TAG[1]));
and5b2 N6P_1_19P_1_I26_1 (.i4(N6P_1_FULL_TAG[1]), .i3(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[3]), .o(N6P_1_CHECK[22]), .i1(N6P_1_FULL_TAG[4]), .i0(N6P_1_FULL_TAG[2]));
and5b2 N6P_1_19P_1_I22_1 (.i4(N6P_1_FULL_TAG[2]), .i3(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[20]), .i1(N6P_1_FULL_TAG[3]), .i0(N6P_1_FULL_TAG[4]));
and5 N6P_1_19P_1_I38_1 (.i4(N6P_1_FULL_TAG[5]), .i2(N6P_1_FULL_TAG[2]), .i3(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[32]), .i0(N6P_1_FULL_TAG[4]), .i1(N6P_1_FULL_TAG[3]));
and5b4 N6P_1_18P_1_I33_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i3(N6P_1_FULL_TAG[2]), .i2(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[1]), .i1(N6P_1_FULL_TAG[4]), .i0(N6P_1_FULL_TAG[3]));
and5b1 N6P_1_18P_1_I39_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i3(N6P_1_FULL_TAG[2]), .i2(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[8]), .i0(N6P_1_FULL_TAG[4]), .i1(N6P_1_FULL_TAG[3]));
and5b1 N6P_1_18P_1_I30_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i3(N6P_1_FULL_TAG[2]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[12]), .i0(N6P_1_FULL_TAG[3]), .i1(N6P_1_FULL_TAG[1]));
and5b1 N6P_1_18P_1_I29_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i3(N6P_1_FULL_TAG[3]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[14]), .i0(N6P_1_FULL_TAG[2]), .i1(N6P_1_FULL_TAG[1]));
and5b1 N6P_1_18P_1_I25_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i3(N6P_1_FULL_TAG[3]), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[15]), .i0(N6P_1_FULL_TAG[1]), .i1(N6P_1_FULL_TAG[2]));
and5b3 N6P_1_18P_1_I37_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[3]), .i3(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[9]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[2]));
and5b3 N6P_1_18P_1_I35_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[4]), .i3(N6P_1_FULL_TAG[3]), .o(N6P_1_CHECK[5]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[2]));
and5b3 N6P_1_18P_1_I34_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[3]), .i3(N6P_1_FULL_TAG[2]), .o(N6P_1_CHECK[3]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[4]));
and5b3 N6P_1_18P_1_I23_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[4]), .i3(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[2]), .i1(N6P_1_FULL_TAG[2]), .i0(N6P_1_FULL_TAG[3]));
and5b2 N6P_1_18P_1_I36_1 (.i4(N6P_1_FULL_TAG[3]), .i3(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[13]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[2]));
and5b2 N6P_1_18P_1_I31_1 (.i4(N6P_1_FULL_TAG[2]), .i3(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[11]), .i1(N6P_1_FULL_TAG[1]), .i0(N6P_1_FULL_TAG[3]));
and5b2 N6P_1_18P_1_I32_1 (.i4(N6P_1_FULL_TAG[1]), .i3(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[4]), .o(N6P_1_CHECK[10]), .i1(N6P_1_FULL_TAG[2]), .i0(N6P_1_FULL_TAG[3]));
and5b2 N6P_1_18P_1_I28_1 (.i4(N6P_1_FULL_TAG[2]), .i3(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[3]), .o(N6P_1_CHECK[7]), .i1(N6P_1_FULL_TAG[4]), .i0(N6P_1_FULL_TAG[1]));
and5b2 N6P_1_18P_1_I26_1 (.i4(N6P_1_FULL_TAG[1]), .i3(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[3]), .o(N6P_1_CHECK[6]), .i1(N6P_1_FULL_TAG[4]), .i0(N6P_1_FULL_TAG[2]));
and5b2 N6P_1_18P_1_I22_1 (.i4(N6P_1_FULL_TAG[2]), .i3(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[4]), .i1(N6P_1_FULL_TAG[3]), .i0(N6P_1_FULL_TAG[4]));
and5 N6P_1_18P_1_I38_1 (.i4(N6P_1_UN_1_D4_16E_18P_E), .i2(N6P_1_FULL_TAG[2]), .i3(N6P_1_FULL_TAG[1]), .o(N6P_1_CHECK[16]), .i0(N6P_1_FULL_TAG[4]), .i1(N6P_1_FULL_TAG[3]));
xor2 N6P_1_17P_1_I34_1_I8_1 (.o(N6P_1_17P_1_I34_1_TQ[0]), .i0(XVDD), .i1(N6P_1_FULL_TAG[0]));
fdce N6P_1_17P_1_I34_1_I7_1 (.d(N6P_1_17P_1_I34_1_TQ[0]), .q(N6P_1_FULL_TAG[0]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND), .gr(RESET_n));
xor2 N6P_1_17P_1_I30_1_I8_1 (.o(N6P_1_17P_1_I30_1_TQ[0]), .i0(N6P_1_17P_1_T4), .i1(N6P_1_FULL_TAG[4]));
fdce N6P_1_17P_1_I30_1_I7_1 (.d(N6P_1_17P_1_I30_1_TQ[0]), .q(N6P_1_FULL_TAG[4]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND), .gr(RESET_n));
xor2 N6P_1_17P_1_I28_1_I8_1 (.o(N6P_1_17P_1_I28_1_TQ[0]), .i0(N6P_1_17P_1_T6), .i1(N6P_1_FULL_TAG[6]));
fdce N6P_1_17P_1_I28_1_I7_1 (.gr(XVDD), .d(N6P_1_17P_1_I28_1_TQ[0]), .q(N6P_1_FULL_TAG[6]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND));
xor2 N6P_1_17P_1_I26_1_I8_1 (.o(N6P_1_17P_1_I26_1_TQ[0]), .i0(N6P_1_FULL_TAG[0]), .i1(N6P_1_FULL_TAG[1]));
fdce N6P_1_17P_1_I26_1_I7_1 (.d(N6P_1_17P_1_I26_1_TQ[0]), .q(N6P_1_FULL_TAG[1]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND), .gr(RESET_n));
xor2 N6P_1_17P_1_I23_1_I8_1 (.o(N6P_1_17P_1_I23_1_TQ[0]), .i0(N6P_1_17P_1_T5), .i1(N6P_1_FULL_TAG[5]));
fdce N6P_1_17P_1_I23_1_I7_1 (.d(N6P_1_17P_1_I23_1_TQ[0]), .q(N6P_1_FULL_TAG[5]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND), .gr(RESET_n));
xor2 N6P_1_17P_1_I20_1_I8_1 (.o(N6P_1_17P_1_I20_1_TQ[0]), .i0(N6P_1_17P_1_T2), .i1(N6P_1_FULL_TAG[2]));
fdce N6P_1_17P_1_I20_1_I7_1 (.d(N6P_1_17P_1_I20_1_TQ[0]), .q(N6P_1_FULL_TAG[2]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND), .gr(RESET_n));
xor2 N6P_1_17P_1_I18_1_I8_1 (.o(N6P_1_17P_1_I18_1_TQ[0]), .i0(N6P_1_17P_1_T3), .i1(N6P_1_FULL_TAG[3]));
fdce N6P_1_17P_1_I18_1_I7_1 (.d(N6P_1_17P_1_I18_1_TQ[0]), .q(N6P_1_FULL_TAG[3]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND), .gr(RESET_n));
xor2 N6P_1_17P_1_I15_1_I8_1 (.o(N6P_1_17P_1_I15_1_TQ[0]), .i0(N6P_1_17P_1_T7), .i1(N6P_1_FULL_TAG[7]));
fdce N6P_1_17P_1_I15_1_I7_1 (.gr(XVDD), .d(N6P_1_17P_1_I15_1_TQ[0]), .q(N6P_1_FULL_TAG[7]), .c(CLK), .ce(UN_1_FD_1_71P_Q), .clr(XGND));
and3 N6P_1_17P_1_I33_1 (.i2(N6P_1_17P_1_T4), .o(N6P_1_17P_1_T6), .i0(N6P_1_FULL_TAG[5]), .i1(N6P_1_FULL_TAG[4]));
and3 N6P_1_17P_1_I32_1 (.i2(N6P_1_FULL_TAG[0]), .o(N6P_1_17P_1_T3), .i0(N6P_1_FULL_TAG[2]), .i1(N6P_1_FULL_TAG[1]));
and5 N6P_1_17P_1_I25_1 (.i4(N6P_1_17P_1_T4), .i2(N6P_1_FULL_TAG[5]), .i3(N6P_1_FULL_TAG[4]), .o(N6P_1_17P_1_TC), .i0(N6P_1_FULL_TAG[7]), .i1(N6P_1_FULL_TAG[6]));
and4 N6P_1_17P_1_I24_1 (.i2(N6P_1_FULL_TAG[4]), .i3(N6P_1_17P_1_T4), .o(N6P_1_17P_1_T7), .i0(N6P_1_FULL_TAG[6]), .i1(N6P_1_FULL_TAG[5]));
and4 N6P_1_17P_1_I16_1 (.i2(N6P_1_FULL_TAG[1]), .i3(N6P_1_FULL_TAG[0]), .o(N6P_1_17P_1_T4), .i0(N6P_1_FULL_TAG[3]), .i1(N6P_1_FULL_TAG[2]));
and2 N6P_1_17P_1_I29_1 (.o(N6P_1_17P_1_T2), .i0(N6P_1_FULL_TAG[1]), .i1(N6P_1_FULL_TAG[0]));
and2 N6P_1_17P_1_I22_1 (.o(N6P_1_17P_1_CEO), .i0(UN_1_FD_1_71P_Q), .i1(N6P_1_17P_1_TC));
and2 N6P_1_17P_1_I21_1 (.o(N6P_1_17P_1_T5), .i0(N6P_1_FULL_TAG[4]), .i1(N6P_1_17P_1_T4));
or4 N6P_1_2P_2 (.i2(N6P_1_UN_2_OR4_2P_I2), .i3(N6P_1_UN_2_OR4_2P_I3), .o(DAV32OR), .i0(N6P_1_UN_2_OR4_2P_I0), .i1(N6P_1_UN_2_OR4_2P_I1));
or4 N6P_1_5P_1 (.i2(N6P_1_UN_1_OR4_5P_I2), .i3(N6P_1_UN_1_OR4_5P_I3), .o(N6P_1_SELECTING), .i0(N6P_1_UN_1_OR4_5P_I0), .i1(N6P_1_UN_1_OR4_5P_I1));
and3b1 N6P_1_60P_1_32 (.i2(N6P_1_CHECK[32]), .o(N6P_1_SELECT[32]), .i0(CHIP_DISABLE[32]), .i1(DAV[32]));
and3b1 N6P_1_60P_1_31 (.i2(DAV[31]), .i0(CHIP_DISABLE[31]), .o(N6P_1_SELECT[31]), .i1(N6P_1_CHECK[31]));
and3b1 N6P_1_60P_1_30 (.i2(DAV[30]), .i0(CHIP_DISABLE[30]), .o(N6P_1_SELECT[30]), .i1(N6P_1_CHECK[30]));
and3b1 N6P_1_60P_1_29 (.i2(DAV[29]), .i0(CHIP_DISABLE[29]), .o(N6P_1_SELECT[29]), .i1(N6P_1_CHECK[29]));
and3b1 N6P_1_60P_1_28 (.i2(DAV[28]), .i0(CHIP_DISABLE[28]), .o(N6P_1_SELECT[28]), .i1(N6P_1_CHECK[28]));
and3b1 N6P_1_60P_1_27 (.i2(DAV[27]), .i0(CHIP_DISABLE[27]), .o(N6P_1_SELECT[27]), .i1(N6P_1_CHECK[27]));
and3b1 N6P_1_60P_1_26 (.i2(DAV[26]), .i0(CHIP_DISABLE[26]), .o(N6P_1_SELECT[26]), .i1(N6P_1_CHECK[26]));
and3b1 N6P_1_60P_1_25 (.i2(DAV[25]), .i0(CHIP_DISABLE[25]), .o(N6P_1_SELECT[25]), .i1(N6P_1_CHECK[25]));
and3b1 N6P_1_60P_1_24 (.i2(DAV[24]), .i0(CHIP_DISABLE[24]), .o(N6P_1_SELECT[24]), .i1(N6P_1_CHECK[24]));
and3b1 N6P_1_60P_1_23 (.i2(DAV[23]), .i0(CHIP_DISABLE[23]), .o(N6P_1_SELECT[23]), .i1(N6P_1_CHECK[23]));
and3b1 N6P_1_60P_1_22 (.i2(DAV[22]), .i0(CHIP_DISABLE[22]), .o(N6P_1_SELECT[22]), .i1(N6P_1_CHECK[22]));
and3b1 N6P_1_60P_1_21 (.i2(DAV[21]), .i0(CHIP_DISABLE[21]), .o(N6P_1_SELECT[21]), .i1(N6P_1_CHECK[21]));
and3b1 N6P_1_60P_1_20 (.i2(DAV[20]), .i0(CHIP_DISABLE[20]), .o(N6P_1_SELECT[20]), .i1(N6P_1_CHECK[20]));
and3b1 N6P_1_60P_1_19 (.i2(DAV[19]), .i0(CHIP_DISABLE[19]), .o(N6P_1_SELECT[19]), .i1(N6P_1_CHECK[19]));
and3b1 N6P_1_60P_1_18 (.i2(DAV[18]), .i0(CHIP_DISABLE[18]), .o(N6P_1_SELECT[18]), .i1(N6P_1_CHECK[18]));
and3b1 N6P_1_60P_1_17 (.i2(DAV[17]), .i0(CHIP_DISABLE[17]), .o(N6P_1_SELECT[17]), .i1(N6P_1_CHECK[17]));
and3b1 N6P_1_60P_1_16 (.i2(DAV[16]), .i0(CHIP_DISABLE[16]), .o(N6P_1_SELECT[16]), .i1(N6P_1_CHECK[16]));
and3b1 N6P_1_60P_1_15 (.i2(DAV[15]), .i0(CHIP_DISABLE[15]), .o(N6P_1_SELECT[15]), .i1(N6P_1_CHECK[15]));
and3b1 N6P_1_60P_1_14 (.i2(DAV[14]), .i0(CHIP_DISABLE[14]), .o(N6P_1_SELECT[14]), .i1(N6P_1_CHECK[14]));
and3b1 N6P_1_60P_1_13 (.i2(DAV[13]), .i0(CHIP_DISABLE[13]), .o(N6P_1_SELECT[13]), .i1(N6P_1_CHECK[13]));
and3b1 N6P_1_60P_1_12 (.i2(DAV[12]), .i0(CHIP_DISABLE[12]), .o(N6P_1_SELECT[12]), .i1(N6P_1_CHECK[12]));
and3b1 N6P_1_60P_1_11 (.i2(DAV[11]), .i0(CHIP_DISABLE[11]), .o(N6P_1_SELECT[11]), .i1(N6P_1_CHECK[11]));
and3b1 N6P_1_60P_1_10 (.i2(DAV[10]), .i0(CHIP_DISABLE[10]), .o(N6P_1_SELECT[10]), .i1(N6P_1_CHECK[10]));
and3b1 N6P_1_60P_1_9 (.i2(DAV[9]), .i0(CHIP_DISABLE[9]), .o(N6P_1_SELECT[9]), .i1(N6P_1_CHECK[9]));
and3b1 N6P_1_60P_1_8 (.i2(DAV[8]), .i0(CHIP_DISABLE[8]), .o(N6P_1_SELECT[8]), .i1(N6P_1_CHECK[8]));
and3b1 N6P_1_60P_1_7 (.i2(DAV[7]), .i0(CHIP_DISABLE[7]), .o(N6P_1_SELECT[7]), .i1(N6P_1_CHECK[7]));
and3b1 N6P_1_60P_1_6 (.i2(DAV[6]), .i0(CHIP_DISABLE[6]), .o(N6P_1_SELECT[6]), .i1(N6P_1_CHECK[6]));
and3b1 N6P_1_60P_1_5 (.i2(DAV[5]), .i0(CHIP_DISABLE[5]), .o(N6P_1_SELECT[5]), .i1(N6P_1_CHECK[5]));
and3b1 N6P_1_60P_1_4 (.i2(DAV[4]), .i0(CHIP_DISABLE[4]), .o(N6P_1_SELECT[4]), .i1(N6P_1_CHECK[4]));
and3b1 N6P_1_60P_1_3 (.i2(DAV[3]), .i0(CHIP_DISABLE[3]), .o(N6P_1_SELECT[3]), .i1(N6P_1_CHECK[3]));
and3b1 N6P_1_60P_1_2 (.i2(DAV[2]), .i0(CHIP_DISABLE[2]), .o(N6P_1_SELECT[2]), .i1(N6P_1_CHECK[2]));
and3b1 N6P_1_60P_1_1 (.i2(DAV[1]), .i0(CHIP_DISABLE[1]), .o(N6P_1_SELECT[1]), .i1(N6P_1_CHECK[1]));
and2 N6P_1_61P_1 (.o(DATA_AVAILABLE), .i0(UN_1_FD_1_71P_Q), .i1(N6P_1_SELECTING));
inv N6P_1_6P_1 (.i(N6P_1_FULL_TAG[5]), .o(N6P_1_UN_1_D4_16E_18P_E));
fdce N66P_1_I8_1_I8_1 (.d(N66P_1_AD), .q(UN_1_BUFG_69P_I), .c(CLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
or3 N66P_1_I12_1 (.i2(N66P_1_A0), .o(N66P_1_AD), .i0(N66P_1_A2), .i1(N66P_1_A1));
and3b2 N66P_1_I10_1 (.i2(UN_1_BUFG_69P_I), .o(N66P_1_A0), .i1(XVDD), .i0(XVDD));
and2b1 N66P_1_I6_1 (.o(N66P_1_A2), .i0(XVDD), .i1(XVDD));
and3b1 N66P_1_I11_1 (.i2(XVDD), .o(N66P_1_A1), .i0(UN_1_BUFG_69P_I), .i1(XVDD));
ifd N77P_1_I6_1 (.d(SQCREG_REQ), .q(CREG_REQ), .c(N77P_1_CB), .gr(RESET_n));
inv N77P_1_I7_1 (.i(CLK), .o(N77P_1_CB));
ifd N64P_1_I6_1_32 (.d(SQDAV[32]), .q(DAV[32]), .c(N64P_1_CB), .gr(RESET_n));
ifd N64P_1_I6_1_31 (.c(N64P_1_CB), .q(DAV[31]), .d(SQDAV[31]), .gr(RESET_n));
ifd N64P_1_I6_1_30 (.c(N64P_1_CB), .q(DAV[30]), .d(SQDAV[30]), .gr(RESET_n));
ifd N64P_1_I6_1_29 (.c(N64P_1_CB), .q(DAV[29]), .d(SQDAV[29]), .gr(RESET_n));
ifd N64P_1_I6_1_28 (.c(N64P_1_CB), .q(DAV[28]), .d(SQDAV[28]), .gr(RESET_n));
ifd N64P_1_I6_1_27 (.c(N64P_1_CB), .q(DAV[27]), .d(SQDAV[27]), .gr(RESET_n));
ifd N64P_1_I6_1_26 (.c(N64P_1_CB), .q(DAV[26]), .d(SQDAV[26]), .gr(RESET_n));
ifd N64P_1_I6_1_25 (.c(N64P_1_CB), .q(DAV[25]), .d(SQDAV[25]), .gr(RESET_n));
ifd N64P_1_I6_1_24 (.c(N64P_1_CB), .q(DAV[24]), .d(SQDAV[24]), .gr(RESET_n));
ifd N64P_1_I6_1_23 (.c(N64P_1_CB), .q(DAV[23]), .d(SQDAV[23]), .gr(RESET_n));
ifd N64P_1_I6_1_22 (.c(N64P_1_CB), .q(DAV[22]), .d(SQDAV[22]), .gr(RESET_n));
ifd N64P_1_I6_1_21 (.c(N64P_1_CB), .q(DAV[21]), .d(SQDAV[21]), .gr(RESET_n));
ifd N64P_1_I6_1_20 (.c(N64P_1_CB), .q(DAV[20]), .d(SQDAV[20]), .gr(RESET_n));
ifd N64P_1_I6_1_19 (.c(N64P_1_CB), .q(DAV[19]), .d(SQDAV[19]), .gr(RESET_n));
ifd N64P_1_I6_1_18 (.c(N64P_1_CB), .q(DAV[18]), .d(SQDAV[18]), .gr(RESET_n));
ifd N64P_1_I6_1_17 (.c(N64P_1_CB), .q(DAV[17]), .d(SQDAV[17]), .gr(RESET_n));
ifd N64P_1_I6_1_16 (.c(N64P_1_CB), .q(DAV[16]), .d(SQDAV[16]), .gr(RESET_n));
ifd N64P_1_I6_1_15 (.c(N64P_1_CB), .q(DAV[15]), .d(SQDAV[15]), .gr(RESET_n));
ifd N64P_1_I6_1_14 (.c(N64P_1_CB), .q(DAV[14]), .d(SQDAV[14]), .gr(RESET_n));
ifd N64P_1_I6_1_13 (.c(N64P_1_CB), .q(DAV[13]), .d(SQDAV[13]), .gr(RESET_n));
ifd N64P_1_I6_1_12 (.c(N64P_1_CB), .q(DAV[12]), .d(SQDAV[12]), .gr(RESET_n));
ifd N64P_1_I6_1_11 (.c(N64P_1_CB), .q(DAV[11]), .d(SQDAV[11]), .gr(RESET_n));
ifd N64P_1_I6_1_10 (.c(N64P_1_CB), .q(DAV[10]), .d(SQDAV[10]), .gr(RESET_n));
ifd N64P_1_I6_1_9 (.c(N64P_1_CB), .q(DAV[9]), .d(SQDAV[9]), .gr(RESET_n));
ifd N64P_1_I6_1_8 (.c(N64P_1_CB), .q(DAV[8]), .d(SQDAV[8]), .gr(RESET_n));
ifd N64P_1_I6_1_7 (.c(N64P_1_CB), .q(DAV[7]), .d(SQDAV[7]), .gr(RESET_n));
ifd N64P_1_I6_1_6 (.c(N64P_1_CB), .q(DAV[6]), .d(SQDAV[6]), .gr(RESET_n));
ifd N64P_1_I6_1_5 (.c(N64P_1_CB), .q(DAV[5]), .d(SQDAV[5]), .gr(RESET_n));
ifd N64P_1_I6_1_4 (.c(N64P_1_CB), .q(DAV[4]), .d(SQDAV[4]), .gr(RESET_n));
ifd N64P_1_I6_1_3 (.c(N64P_1_CB), .q(DAV[3]), .d(SQDAV[3]), .gr(RESET_n));
ifd N64P_1_I6_1_2 (.c(N64P_1_CB), .q(DAV[2]), .d(SQDAV[2]), .gr(RESET_n));
ifd N64P_1_I6_1_1 (.c(N64P_1_CB), .q(DAV[1]), .d(SQDAV[1]), .gr(RESET_n));
inv N64P_1_I7_1 (.i(CLKD2), .o(N64P_1_CB));
fdce N47P_1_15P_1_I4_1_32 (.d(N47P_1_DIN[31]), .q(CHIP_DISABLE[32]), .c(N47P_1_15P_1_CB), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_31 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[31]), .d(N47P_1_DIN[30]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_30 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[30]), .d(N47P_1_DIN[29]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_29 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[29]), .d(N47P_1_DIN[28]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_28 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[28]), .d(N47P_1_DIN[27]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_27 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[27]), .d(N47P_1_DIN[26]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_26 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[26]), .d(N47P_1_DIN[25]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_25 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[25]), .d(N47P_1_DIN[24]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_24 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[24]), .d(N47P_1_DIN[23]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_23 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[23]), .d(N47P_1_DIN[22]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_22 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[22]), .d(N47P_1_DIN[21]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_21 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[21]), .d(N47P_1_DIN[20]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_20 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[20]), .d(N47P_1_DIN[19]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_19 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[19]), .d(N47P_1_DIN[18]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_18 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[18]), .d(N47P_1_DIN[17]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_17 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[17]), .d(N47P_1_DIN[16]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_16 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[16]), .d(N47P_1_DIN[15]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_15 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[15]), .d(N47P_1_DIN[14]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_14 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[14]), .d(N47P_1_DIN[13]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_13 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[13]), .d(N47P_1_DIN[12]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_12 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[12]), .d(N47P_1_DIN[11]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_11 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[11]), .d(N47P_1_DIN[10]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_10 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[10]), .d(N47P_1_DIN[9]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_9 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[9]), .d(N47P_1_DIN[8]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_8 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[8]), .d(N47P_1_DIN[7]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_7 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[7]), .d(N47P_1_DIN[6]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_6 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[6]), .d(N47P_1_DIN[5]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_5 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[5]), .d(N47P_1_DIN[4]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_4 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[4]), .d(N47P_1_DIN[3]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_3 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[3]), .d(N47P_1_DIN[2]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_2 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[2]), .d(N47P_1_DIN[1]), .gr(RESET_n));
fdce N47P_1_15P_1_I4_1_1 (.clr(XGND), .ce(XVDD), .c(N47P_1_15P_1_CB), .q(CHIP_DISABLE[1]), .d(N47P_1_DIN[0]), .gr(RESET_n));
inv N47P_1_15P_1_I5_1 (.i(N47P_1_REG_CDIS_WR_n), .o(N47P_1_15P_1_CB));
inv N47P_1_16P_1_21P_1 (.i(N47P_1_16P_1_UN_1_INV_21P_I), .o(N47P_1_16P_1_UN_1_INV_20P_I));
inv N47P_1_16P_1_22P_1 (.i(N47P_1_UN_1_DELAY_16P_DELAY), .o(N47P_1_16P_1_UN_1_INV_21P_I));
inv N47P_1_16P_1_20P_1 (.i(N47P_1_16P_1_UN_1_INV_20P_I), .o(N47P_1_16P_1_UN_1_INV_14P_I));
inv N47P_1_16P_1_19P_1 (.i(N47P_1_16P_1_UN_1_INV_18P_O), .o(N47P_1_16P_1_UN_1_INV_13P_I));
inv N47P_1_16P_1_18P_1 (.i(N47P_1_16P_1_UN_1_INV_17P_O), .o(N47P_1_16P_1_UN_1_INV_18P_O));
inv N47P_1_16P_1_17P_1 (.i(N47P_1_16P_1_UN_1_INV_16P_O), .o(N47P_1_16P_1_UN_1_INV_17P_O));
inv N47P_1_16P_1_16P_1 (.i(N47P_1_16P_1_UN_1_INV_15P_O), .o(N47P_1_16P_1_UN_1_INV_16P_O));
inv N47P_1_16P_1_15P_1 (.i(N47P_1_16P_1_UN_1_INV_14P_O), .o(N47P_1_16P_1_UN_1_INV_15P_O));
inv N47P_1_16P_1_14P_1 (.i(N47P_1_16P_1_UN_1_INV_14P_I), .o(N47P_1_16P_1_UN_1_INV_14P_O));
inv N47P_1_16P_1_13P_1 (.i(N47P_1_16P_1_UN_1_INV_13P_I), .o(N47P_1_REG_CDIS_WR_n));
obuft N47P_1_3P_1_32 (.i(N47P_1_DOUT[31]), .o(SQD[31]), .t(REG_RD_n));
obuft N47P_1_3P_1_31 (.t(REG_RD_n), .o(SQD[30]), .i(N47P_1_DOUT[30]));
obuft N47P_1_3P_1_30 (.t(REG_RD_n), .o(SQD[29]), .i(N47P_1_DOUT[29]));
obuft N47P_1_3P_1_29 (.t(REG_RD_n), .o(SQD[28]), .i(N47P_1_DOUT[28]));
obuft N47P_1_3P_1_28 (.t(REG_RD_n), .o(SQD[27]), .i(N47P_1_DOUT[27]));
obuft N47P_1_3P_1_27 (.t(REG_RD_n), .o(SQD[26]), .i(N47P_1_DOUT[26]));
obuft N47P_1_3P_1_26 (.t(REG_RD_n), .o(SQD[25]), .i(N47P_1_DOUT[25]));
obuft N47P_1_3P_1_25 (.t(REG_RD_n), .o(SQD[24]), .i(N47P_1_DOUT[24]));
obuft N47P_1_3P_1_24 (.t(REG_RD_n), .o(SQD[23]), .i(N47P_1_DOUT[23]));
obuft N47P_1_3P_1_23 (.t(REG_RD_n), .o(SQD[22]), .i(N47P_1_DOUT[22]));
obuft N47P_1_3P_1_22 (.t(REG_RD_n), .o(SQD[21]), .i(N47P_1_DOUT[21]));
obuft N47P_1_3P_1_21 (.t(REG_RD_n), .o(SQD[20]), .i(N47P_1_DOUT[20]));
obuft N47P_1_3P_1_20 (.t(REG_RD_n), .o(SQD[19]), .i(N47P_1_DOUT[19]));
obuft N47P_1_3P_1_19 (.t(REG_RD_n), .o(SQD[18]), .i(N47P_1_DOUT[18]));
obuft N47P_1_3P_1_18 (.t(REG_RD_n), .o(SQD[17]), .i(N47P_1_DOUT[17]));
obuft N47P_1_3P_1_17 (.t(REG_RD_n), .o(SQD[16]), .i(N47P_1_DOUT[16]));
obuft N47P_1_3P_1_16 (.t(REG_RD_n), .o(SQD[15]), .i(N47P_1_DOUT[15]));
obuft N47P_1_3P_1_15 (.t(REG_RD_n), .o(SQD[14]), .i(N47P_1_DOUT[14]));
obuft N47P_1_3P_1_14 (.t(REG_RD_n), .o(SQD[13]), .i(N47P_1_DOUT[13]));
obuft N47P_1_3P_1_13 (.t(REG_RD_n), .o(SQD[12]), .i(N47P_1_DOUT[12]));
obuft N47P_1_3P_1_12 (.t(REG_RD_n), .o(SQD[11]), .i(N47P_1_DOUT[11]));
obuft N47P_1_3P_1_11 (.t(REG_RD_n), .o(SQD[10]), .i(N47P_1_DOUT[10]));
obuft N47P_1_3P_1_10 (.t(REG_RD_n), .o(SQD[9]), .i(N47P_1_DOUT[9]));
obuft N47P_1_3P_1_9 (.t(REG_RD_n), .o(SQD[8]), .i(N47P_1_DOUT[8]));
obuft N47P_1_3P_1_8 (.t(REG_RD_n), .o(SQD[7]), .i(N47P_1_DOUT[7]));
obuft N47P_1_3P_1_7 (.t(REG_RD_n), .o(SQD[6]), .i(N47P_1_DOUT[6]));
obuft N47P_1_3P_1_6 (.t(REG_RD_n), .o(SQD[5]), .i(N47P_1_DOUT[5]));
obuft N47P_1_3P_1_5 (.t(REG_RD_n), .o(SQD[4]), .i(N47P_1_DOUT[4]));
obuft N47P_1_3P_1_4 (.t(REG_RD_n), .o(SQD[3]), .i(N47P_1_DOUT[3]));
obuft N47P_1_3P_1_3 (.t(REG_RD_n), .o(SQD[2]), .i(N47P_1_DOUT[2]));
obuft N47P_1_3P_1_2 (.t(REG_RD_n), .o(SQD[1]), .i(N47P_1_DOUT[1]));
obuft N47P_1_3P_1_1 (.t(REG_RD_n), .o(SQD[0]), .i(N47P_1_DOUT[0]));
and4b3 N47P_1_12P_1 (.i2(REG_SEL[1]), .i3(REG_SEL[2]), .o(N47P_1_CDIS_REG_RD), .i1(REG_RD_n), .i0(REG_SEL[0]));
nand4b3 N47P_1_14P_1 (.i2(REG_SEL[1]), .i3(REG_SEL[2]), .o(N47P_1_UN_1_DELAY_16P_DELAY), .i1(REG_WR_n), .i0(REG_SEL[0]));
and2 N47P_1_11P_1_32 (.o(N47P_1_DOUT[31]), .i0(N47P_1_CDIS_REG_RD), .i1(CHIP_DISABLE[32]));
and2 N47P_1_11P_1_31 (.i1(CHIP_DISABLE[31]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[30]));
and2 N47P_1_11P_1_30 (.i1(CHIP_DISABLE[30]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[29]));
and2 N47P_1_11P_1_29 (.i1(CHIP_DISABLE[29]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[28]));
and2 N47P_1_11P_1_28 (.i1(CHIP_DISABLE[28]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[27]));
and2 N47P_1_11P_1_27 (.i1(CHIP_DISABLE[27]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[26]));
and2 N47P_1_11P_1_26 (.i1(CHIP_DISABLE[26]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[25]));
and2 N47P_1_11P_1_25 (.i1(CHIP_DISABLE[25]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[24]));
and2 N47P_1_11P_1_24 (.i1(CHIP_DISABLE[24]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[23]));
and2 N47P_1_11P_1_23 (.i1(CHIP_DISABLE[23]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[22]));
and2 N47P_1_11P_1_22 (.i1(CHIP_DISABLE[22]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[21]));
and2 N47P_1_11P_1_21 (.i1(CHIP_DISABLE[21]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[20]));
and2 N47P_1_11P_1_20 (.i1(CHIP_DISABLE[20]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[19]));
and2 N47P_1_11P_1_19 (.i1(CHIP_DISABLE[19]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[18]));
and2 N47P_1_11P_1_18 (.i1(CHIP_DISABLE[18]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[17]));
and2 N47P_1_11P_1_17 (.i1(CHIP_DISABLE[17]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[16]));
and2 N47P_1_11P_1_16 (.i1(CHIP_DISABLE[16]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[15]));
and2 N47P_1_11P_1_15 (.i1(CHIP_DISABLE[15]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[14]));
and2 N47P_1_11P_1_14 (.i1(CHIP_DISABLE[14]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[13]));
and2 N47P_1_11P_1_13 (.i1(CHIP_DISABLE[13]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[12]));
and2 N47P_1_11P_1_12 (.i1(CHIP_DISABLE[12]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[11]));
and2 N47P_1_11P_1_11 (.i1(CHIP_DISABLE[11]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[10]));
and2 N47P_1_11P_1_10 (.i1(CHIP_DISABLE[10]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[9]));
and2 N47P_1_11P_1_9 (.i1(CHIP_DISABLE[9]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[8]));
and2 N47P_1_11P_1_8 (.i1(CHIP_DISABLE[8]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[7]));
and2 N47P_1_11P_1_7 (.i1(CHIP_DISABLE[7]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[6]));
and2 N47P_1_11P_1_6 (.i1(CHIP_DISABLE[6]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[5]));
and2 N47P_1_11P_1_5 (.i1(CHIP_DISABLE[5]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[4]));
and2 N47P_1_11P_1_4 (.i1(CHIP_DISABLE[4]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[3]));
and2 N47P_1_11P_1_3 (.i1(CHIP_DISABLE[3]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[2]));
and2 N47P_1_11P_1_2 (.i1(CHIP_DISABLE[2]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[1]));
and2 N47P_1_11P_1_1 (.i1(CHIP_DISABLE[1]), .i0(N47P_1_CDIS_REG_RD), .o(N47P_1_DOUT[0]));
ibuf N47P_1_2P_1_32 (.i(SQD[31]), .o(N47P_1_DIN[31]));
ibuf N47P_1_2P_1_31 (.o(N47P_1_DIN[30]), .i(SQD[30]));
ibuf N47P_1_2P_1_30 (.o(N47P_1_DIN[29]), .i(SQD[29]));
ibuf N47P_1_2P_1_29 (.o(N47P_1_DIN[28]), .i(SQD[28]));
ibuf N47P_1_2P_1_28 (.o(N47P_1_DIN[27]), .i(SQD[27]));
ibuf N47P_1_2P_1_27 (.o(N47P_1_DIN[26]), .i(SQD[26]));
ibuf N47P_1_2P_1_26 (.o(N47P_1_DIN[25]), .i(SQD[25]));
ibuf N47P_1_2P_1_25 (.o(N47P_1_DIN[24]), .i(SQD[24]));
ibuf N47P_1_2P_1_24 (.o(N47P_1_DIN[23]), .i(SQD[23]));
ibuf N47P_1_2P_1_23 (.o(N47P_1_DIN[22]), .i(SQD[22]));
ibuf N47P_1_2P_1_22 (.o(N47P_1_DIN[21]), .i(SQD[21]));
ibuf N47P_1_2P_1_21 (.o(N47P_1_DIN[20]), .i(SQD[20]));
ibuf N47P_1_2P_1_20 (.o(N47P_1_DIN[19]), .i(SQD[19]));
ibuf N47P_1_2P_1_19 (.o(N47P_1_DIN[18]), .i(SQD[18]));
ibuf N47P_1_2P_1_18 (.o(N47P_1_DIN[17]), .i(SQD[17]));
ibuf N47P_1_2P_1_17 (.o(N47P_1_DIN[16]), .i(SQD[16]));
ibuf N47P_1_2P_1_16 (.o(N47P_1_DIN[15]), .i(SQD[15]));
ibuf N47P_1_2P_1_15 (.o(N47P_1_DIN[14]), .i(SQD[14]));
ibuf N47P_1_2P_1_14 (.o(N47P_1_DIN[13]), .i(SQD[13]));
ibuf N47P_1_2P_1_13 (.o(N47P_1_DIN[12]), .i(SQD[12]));
ibuf N47P_1_2P_1_12 (.o(N47P_1_DIN[11]), .i(SQD[11]));
ibuf N47P_1_2P_1_11 (.o(N47P_1_DIN[10]), .i(SQD[10]));
ibuf N47P_1_2P_1_10 (.o(N47P_1_DIN[9]), .i(SQD[9]));
ibuf N47P_1_2P_1_9 (.o(N47P_1_DIN[8]), .i(SQD[8]));
ibuf N47P_1_2P_1_8 (.o(N47P_1_DIN[7]), .i(SQD[7]));
ibuf N47P_1_2P_1_7 (.o(N47P_1_DIN[6]), .i(SQD[6]));
ibuf N47P_1_2P_1_6 (.o(N47P_1_DIN[5]), .i(SQD[5]));
ibuf N47P_1_2P_1_5 (.o(N47P_1_DIN[4]), .i(SQD[4]));
ibuf N47P_1_2P_1_4 (.o(N47P_1_DIN[3]), .i(SQD[3]));
ibuf N47P_1_2P_1_3 (.o(N47P_1_DIN[2]), .i(SQD[2]));
ibuf N47P_1_2P_1_2 (.o(N47P_1_DIN[1]), .i(SQD[1]));
ibuf N47P_1_2P_1_1 (.o(N47P_1_DIN[0]), .i(SQD[0]));
fdce N31P_1_4P_1_19P_1_I14_1_I7_1_I7_1_I6_1 (.gr(XVDD), .d(N31P_1_4P_1_19P_1_I14_1_I7_1_QD[0]), .q(N31P_1_4P_1_S[3]), .c(CLK), .ce(XVDD), .clr(XGND));
or2 N31P_1_4P_1_19P_1_I14_1_I7_1_I9_1 (.o(N31P_1_4P_1_19P_1_I14_1_I7_1_QD[0]), .i0(N31P_1_4P_1_19P_1_I14_1_I7_1_A1[0]), .i1(N31P_1_4P_1_19P_1_I14_1_I7_1_A0));
and3b2 N31P_1_4P_1_19P_1_I14_1_I7_1_I8_1 (.i2(N31P_1_4P_1_S[3]), .o(N31P_1_4P_1_19P_1_I14_1_I7_1_A0), .i1(N31P_1_4P_1_19P_1_I14_1_CE_S), .i0(XGND));
and3b1 N31P_1_4P_1_19P_1_I14_1_I7_1_I10_1 (.i2(N31P_1_4P_1_19P_1_I14_1_CE_S), .o(N31P_1_4P_1_19P_1_I14_1_I7_1_A1[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I14_1_D_S[0]));
xor2 N31P_1_4P_1_19P_1_I14_1_I9_1 (.o(N31P_1_4P_1_19P_1_I14_1_TQ), .i0(N31P_1_4P_1_19P_1_T3), .i1(N31P_1_4P_1_S[3]));
or2 N31P_1_4P_1_19P_1_I14_1_I12_1 (.o(N31P_1_4P_1_19P_1_I14_1_CE_S), .i0(N31P_1_4P_1_CLK_ENA), .i1(XGND));
or2 N31P_1_4P_1_19P_1_I14_1_I11_1 (.o(N31P_1_4P_1_19P_1_I14_1_D_S[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I14_1_TQ));
fdce N31P_1_4P_1_19P_1_I13_1_I7_1_I7_1_I6_1 (.d(N31P_1_4P_1_19P_1_I13_1_I7_1_QD[0]), .q(N31P_1_4P_1_S[0]), .c(CLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
or2 N31P_1_4P_1_19P_1_I13_1_I7_1_I9_1 (.o(N31P_1_4P_1_19P_1_I13_1_I7_1_QD[0]), .i0(N31P_1_4P_1_19P_1_I13_1_I7_1_A1[0]), .i1(N31P_1_4P_1_19P_1_I13_1_I7_1_A0));
and3b2 N31P_1_4P_1_19P_1_I13_1_I7_1_I8_1 (.i2(N31P_1_4P_1_S[0]), .o(N31P_1_4P_1_19P_1_I13_1_I7_1_A0), .i1(N31P_1_4P_1_19P_1_I13_1_CE_S), .i0(XGND));
and3b1 N31P_1_4P_1_19P_1_I13_1_I7_1_I10_1 (.i2(N31P_1_4P_1_19P_1_I13_1_CE_S), .o(N31P_1_4P_1_19P_1_I13_1_I7_1_A1[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I13_1_D_S[0]));
xor2 N31P_1_4P_1_19P_1_I13_1_I9_1 (.o(N31P_1_4P_1_19P_1_I13_1_TQ), .i0(XVDD), .i1(N31P_1_4P_1_S[0]));
or2 N31P_1_4P_1_19P_1_I13_1_I12_1 (.o(N31P_1_4P_1_19P_1_I13_1_CE_S), .i0(N31P_1_4P_1_CLK_ENA), .i1(XGND));
or2 N31P_1_4P_1_19P_1_I13_1_I11_1 (.o(N31P_1_4P_1_19P_1_I13_1_D_S[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I13_1_TQ));
fdce N31P_1_4P_1_19P_1_I18_1_I7_1_I7_1_I6_1 (.d(N31P_1_4P_1_19P_1_I18_1_I7_1_QD[0]), .q(N31P_1_4P_1_S[1]), .c(CLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
or2 N31P_1_4P_1_19P_1_I18_1_I7_1_I9_1 (.o(N31P_1_4P_1_19P_1_I18_1_I7_1_QD[0]), .i0(N31P_1_4P_1_19P_1_I18_1_I7_1_A1[0]), .i1(N31P_1_4P_1_19P_1_I18_1_I7_1_A0));
and3b2 N31P_1_4P_1_19P_1_I18_1_I7_1_I8_1 (.i2(N31P_1_4P_1_S[1]), .o(N31P_1_4P_1_19P_1_I18_1_I7_1_A0), .i1(N31P_1_4P_1_19P_1_I18_1_CE_S), .i0(XGND));
and3b1 N31P_1_4P_1_19P_1_I18_1_I7_1_I10_1 (.i2(N31P_1_4P_1_19P_1_I18_1_CE_S), .o(N31P_1_4P_1_19P_1_I18_1_I7_1_A1[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I18_1_D_S[0]));
xor2 N31P_1_4P_1_19P_1_I18_1_I9_1 (.o(N31P_1_4P_1_19P_1_I18_1_TQ), .i0(N31P_1_4P_1_S[0]), .i1(N31P_1_4P_1_S[1]));
or2 N31P_1_4P_1_19P_1_I18_1_I12_1 (.o(N31P_1_4P_1_19P_1_I18_1_CE_S), .i0(N31P_1_4P_1_CLK_ENA), .i1(XGND));
or2 N31P_1_4P_1_19P_1_I18_1_I11_1 (.o(N31P_1_4P_1_19P_1_I18_1_D_S[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I18_1_TQ));
fdce N31P_1_4P_1_19P_1_I15_1_I7_1_I7_1_I6_1 (.d(N31P_1_4P_1_19P_1_I15_1_I7_1_QD[0]), .q(N31P_1_4P_1_S[2]), .c(CLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
or2 N31P_1_4P_1_19P_1_I15_1_I7_1_I9_1 (.o(N31P_1_4P_1_19P_1_I15_1_I7_1_QD[0]), .i0(N31P_1_4P_1_19P_1_I15_1_I7_1_A1[0]), .i1(N31P_1_4P_1_19P_1_I15_1_I7_1_A0));
and3b2 N31P_1_4P_1_19P_1_I15_1_I7_1_I8_1 (.i2(N31P_1_4P_1_S[2]), .o(N31P_1_4P_1_19P_1_I15_1_I7_1_A0), .i1(N31P_1_4P_1_19P_1_I15_1_CE_S), .i0(XGND));
and3b1 N31P_1_4P_1_19P_1_I15_1_I7_1_I10_1 (.i2(N31P_1_4P_1_19P_1_I15_1_CE_S), .o(N31P_1_4P_1_19P_1_I15_1_I7_1_A1[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I15_1_D_S[0]));
xor2 N31P_1_4P_1_19P_1_I15_1_I9_1 (.o(N31P_1_4P_1_19P_1_I15_1_TQ), .i0(N31P_1_4P_1_19P_1_T2), .i1(N31P_1_4P_1_S[2]));
or2 N31P_1_4P_1_19P_1_I15_1_I12_1 (.o(N31P_1_4P_1_19P_1_I15_1_CE_S), .i0(N31P_1_4P_1_CLK_ENA), .i1(XGND));
or2 N31P_1_4P_1_19P_1_I15_1_I11_1 (.o(N31P_1_4P_1_19P_1_I15_1_D_S[0]), .i0(XGND), .i1(N31P_1_4P_1_19P_1_I15_1_TQ));
and3 N31P_1_4P_1_19P_1_I11_1 (.i2(N31P_1_4P_1_S[0]), .o(N31P_1_4P_1_19P_1_T3), .i0(N31P_1_4P_1_S[2]), .i1(N31P_1_4P_1_S[1]));
and4 N31P_1_4P_1_19P_1_I16_1 (.i2(N31P_1_4P_1_S[1]), .i3(N31P_1_4P_1_S[0]), .o(N31P_1_4P_1_19P_1_TC), .i0(N31P_1_4P_1_S[3]), .i1(N31P_1_4P_1_S[2]));
and2 N31P_1_4P_1_19P_1_I17_1 (.o(N31P_1_4P_1_19P_1_T2), .i0(N31P_1_4P_1_S[1]), .i1(N31P_1_4P_1_S[0]));
and2 N31P_1_4P_1_19P_1_I10_1 (.o(N31P_1_4P_1_19P_1_CEO), .i0(N31P_1_4P_1_CLK_ENA), .i1(N31P_1_4P_1_19P_1_TC));
and4b2 N31P_1_4P_1_23P_1_I17_1 (.i3(N31P_1_4P_1_S[1]), .i2(XVDD), .o(N31P_1_4P_1_C[0]), .i1(N31P_1_4P_1_S[2]), .i0(N31P_1_4P_1_S[0]));
and4b2 N31P_1_4P_1_23P_1_I14_1 (.i3(N31P_1_4P_1_S[0]), .i2(XVDD), .o(N31P_1_4P_1_STAGE[1]), .i1(N31P_1_4P_1_S[2]), .i0(N31P_1_4P_1_S[1]));
and4b2 N31P_1_4P_1_23P_1_I18_1 (.i3(N31P_1_4P_1_S[2]), .i2(XVDD), .o(N31P_1_4P_1_STAGE[2]), .i1(N31P_1_4P_1_S[1]), .i0(N31P_1_4P_1_S[0]));
and4b1 N31P_1_4P_1_23P_1_I13_1 (.i3(N31P_1_4P_1_S[1]), .i2(XVDD), .o(N31P_1_4P_1_C[3]), .i0(N31P_1_4P_1_S[0]), .i1(N31P_1_4P_1_S[2]));
and4b1 N31P_1_4P_1_23P_1_I16_1 (.i3(N31P_1_4P_1_S[1]), .i2(XVDD), .o(N31P_1_4P_1_C[1]), .i0(N31P_1_4P_1_S[2]), .i1(N31P_1_4P_1_S[0]));
and4b1 N31P_1_4P_1_23P_1_I15_1 (.i3(N31P_1_4P_1_S[0]), .i2(XVDD), .o(N31P_1_4P_1_C[2]), .i0(N31P_1_4P_1_S[1]), .i1(N31P_1_4P_1_S[2]));
and4 N31P_1_4P_1_23P_1_I22_1 (.i2(N31P_1_4P_1_S[0]), .i3(XVDD), .o(N31P_1_4P_1_STAGE[3]), .i0(N31P_1_4P_1_S[2]), .i1(N31P_1_4P_1_S[1]));
and4b3 N31P_1_4P_1_23P_1_I23_1 (.i2(N31P_1_4P_1_S[0]), .i3(XVDD), .o(N31P_1_ALL_DATA_PROCESSED), .i1(N31P_1_4P_1_S[2]), .i0(N31P_1_4P_1_S[1]));
fdce N31P_1_4P_1_32P_1_I8_1 (.d(XVDD), .q(N31P_1_4P_1_UN_1_FDC_32P_Q), .c(N31P_1_DATA_READY), .ce(XVDD), .clr(N31P_1_4P_1_STAGE[1]), .gr(RESET_n));
or5 N31P_1_4P_1_31P_1 (.i4(N31P_1_4P_1_UN_1_FDC_32P_Q), .i2(N31P_1_4P_1_C[2]), .i3(N31P_1_4P_1_C[3]), .o(N31P_1_4P_1_UN_1_OR4_30P_I3), .i0(N31P_1_4P_1_C[0]), .i1(N31P_1_4P_1_C[1]));
and3 N31P_1_4P_1_20P_1 (.i2(ENW_[1]), .o(MEMORY_REQUEST_n), .i0(ENW_[3]), .i1(ENW_[2]));
or4 N31P_1_4P_1_30P_1 (.i2(N31P_1_4P_1_UN_1_AND2B1_29P_O), .i3(N31P_1_4P_1_UN_1_OR4_30P_I3), .o(N31P_1_4P_1_CLK_ENA), .i0(N31P_1_4P_1_UN_1_AND2B1_27P_O), .i1(N31P_1_4P_1_UN_1_AND2B1_28P_O));
and2b1 N31P_1_4P_1_27P_1 (.o(N31P_1_4P_1_UN_1_AND2B1_27P_O), .i0(MEMORY_ACK_n), .i1(N31P_1_4P_1_STAGE[3]));
and2b1 N31P_1_4P_1_29P_1 (.o(N31P_1_4P_1_UN_1_AND2B1_29P_O), .i0(MEMORY_ACK_n), .i1(N31P_1_4P_1_STAGE[1]));
and2b1 N31P_1_4P_1_28P_1 (.o(N31P_1_4P_1_UN_1_AND2B1_28P_O), .i0(MEMORY_ACK_n), .i1(N31P_1_4P_1_STAGE[2]));
inv N31P_1_4P_1_5P_1 (.i(N31P_1_4P_1_STAGE[1]), .o(ENW_[1]));
inv N31P_1_4P_1_4P_1 (.i(N31P_1_4P_1_STAGE[2]), .o(ENW_[2]));
inv N31P_1_4P_1_3P_1 (.i(N31P_1_4P_1_STAGE[3]), .o(ENW_[3]));
fdce N31P_1_42P_1_I8_1 (.d(XVDD), .q(N31P_1_UN_1_FDC_42P_Q), .c(CREG_REQ), .ce(XVDD), .clr(LATCH[4]), .gr(RESET_n));
fdce N31P_1_40P_1_I8_1 (.d(LATCH_TAG), .q(CADD_ENABLE), .c(CREG_REQ), .ce(XVDD), .clr(N31P_1_CMOS_END), .gr(RESET_n));
and4b2 N31P_1_2P_1_52P_1_I17_1 (.i3(N31P_1_2P_1_STATES[2]), .i2(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(N31P_1_2P_1_WAIT[1]), .i1(N31P_1_2P_1_STATES[3]), .i0(N31P_1_2P_1_STATES[1]));
and4b2 N31P_1_2P_1_52P_1_I14_1 (.i3(N31P_1_2P_1_STATES[1]), .i2(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(N31P_1_2P_1_WAIT[0]), .i1(N31P_1_2P_1_STATES[3]), .i0(N31P_1_2P_1_STATES[2]));
and4b2 N31P_1_2P_1_52P_1_I18_1 (.i3(N31P_1_2P_1_STATES[3]), .i2(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(N31P_1_2P_1_WAIT[3]), .i1(N31P_1_2P_1_STATES[2]), .i0(N31P_1_2P_1_STATES[1]));
and4b1 N31P_1_2P_1_52P_1_I13_1 (.i3(N31P_1_2P_1_STATES[2]), .i2(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(N31P_1_2P_1_WAIT[4]), .i0(N31P_1_2P_1_STATES[1]), .i1(N31P_1_2P_1_STATES[3]));
and4b1 N31P_1_2P_1_52P_1_I16_1 (.i3(N31P_1_2P_1_STATES[2]), .i2(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(N31P_1_2P_1_WAIT[2]), .i0(N31P_1_2P_1_STATES[3]), .i1(N31P_1_2P_1_STATES[1]));
and4b1 N31P_1_2P_1_52P_1_I15_1 (.i3(N31P_1_2P_1_STATES[1]), .i2(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(CONVERT_START), .i0(N31P_1_2P_1_STATES[2]), .i1(N31P_1_2P_1_STATES[3]));
and4 N31P_1_2P_1_52P_1_I22_1 (.i2(N31P_1_2P_1_STATES[1]), .i3(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(N31P_1_2P_1_WAIT[5]), .i0(N31P_1_2P_1_STATES[3]), .i1(N31P_1_2P_1_STATES[2]));
and4b3 N31P_1_2P_1_52P_1_I23_1 (.i2(N31P_1_2P_1_STATES[1]), .i3(N31P_1_2P_1_UN_1_D3_8E_52P_E), .o(LATCH_TAG), .i1(N31P_1_2P_1_STATES[3]), .i0(N31P_1_2P_1_STATES[2]));
and4b2 N31P_1_2P_1_51P_1_I17_1 (.i3(N31P_1_2P_1_STATES[2]), .i2(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(N31P_1_2P_1_STROBE[2]), .i1(N31P_1_2P_1_STATES[3]), .i0(N31P_1_2P_1_STATES[1]));
and4b2 N31P_1_2P_1_51P_1_I14_1 (.i3(N31P_1_2P_1_STATES[1]), .i2(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(LATCH[1]), .i1(N31P_1_2P_1_STATES[3]), .i0(N31P_1_2P_1_STATES[2]));
and4b2 N31P_1_2P_1_51P_1_I18_1 (.i3(N31P_1_2P_1_STATES[3]), .i2(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(N31P_1_2P_1_STROBE[3]), .i1(N31P_1_2P_1_STATES[2]), .i0(N31P_1_2P_1_STATES[1]));
and4b1 N31P_1_2P_1_51P_1_I13_1 (.i3(N31P_1_2P_1_STATES[2]), .i2(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(N31P_1_2P_1_STROBE[4]), .i0(N31P_1_2P_1_STATES[1]), .i1(N31P_1_2P_1_STATES[3]));
and4b1 N31P_1_2P_1_51P_1_I16_1 (.i3(N31P_1_2P_1_STATES[2]), .i2(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(LATCH[2]), .i0(N31P_1_2P_1_STATES[3]), .i1(N31P_1_2P_1_STATES[1]));
and4b1 N31P_1_2P_1_51P_1_I15_1 (.i3(N31P_1_2P_1_STATES[1]), .i2(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(LATCH[3]), .i0(N31P_1_2P_1_STATES[2]), .i1(N31P_1_2P_1_STATES[3]));
and4 N31P_1_2P_1_51P_1_I22_1 (.i2(N31P_1_2P_1_STATES[1]), .i3(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(LATCH[4]), .i0(N31P_1_2P_1_STATES[3]), .i1(N31P_1_2P_1_STATES[2]));
and4b3 N31P_1_2P_1_51P_1_I23_1 (.i2(N31P_1_2P_1_STATES[1]), .i3(N31P_1_2P_1_UN_1_D3_8E_51P_E), .o(N31P_1_2P_1_STROBE[1]), .i1(N31P_1_2P_1_STATES[3]), .i0(N31P_1_2P_1_STATES[2]));
xor2 N31P_1_2P_1_83P_1_I34_1_I8_1 (.o(N31P_1_2P_1_83P_1_I34_1_TQ[0]), .i0(XVDD), .i1(N31P_1_2P_1_STATES[0]));
fdce N31P_1_2P_1_83P_1_I34_1_I7_1 (.d(N31P_1_2P_1_83P_1_I34_1_TQ[0]), .q(N31P_1_2P_1_STATES[0]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE), .gr(RESET_n));
xor2 N31P_1_2P_1_83P_1_I30_1_I8_1 (.o(N31P_1_2P_1_83P_1_I30_1_TQ[0]), .i0(N31P_1_2P_1_83P_1_T4), .i1(N31P_1_2P_1_STATES[4]));
fdce N31P_1_2P_1_83P_1_I30_1_I7_1 (.d(N31P_1_2P_1_83P_1_I30_1_TQ[0]), .q(N31P_1_2P_1_STATES[4]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE), .gr(RESET_n));
xor2 N31P_1_2P_1_83P_1_I28_1_I8_1 (.o(N31P_1_2P_1_83P_1_I28_1_TQ[0]), .i0(N31P_1_2P_1_83P_1_T6), .i1(N31P_1_2P_1_STATES[6]));
fdce N31P_1_2P_1_83P_1_I28_1_I7_1 (.gr(XVDD), .d(N31P_1_2P_1_83P_1_I28_1_TQ[0]), .q(N31P_1_2P_1_STATES[6]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE));
xor2 N31P_1_2P_1_83P_1_I26_1_I8_1 (.o(N31P_1_2P_1_83P_1_I26_1_TQ[0]), .i0(N31P_1_2P_1_STATES[0]), .i1(N31P_1_2P_1_STATES[1]));
fdce N31P_1_2P_1_83P_1_I26_1_I7_1 (.d(N31P_1_2P_1_83P_1_I26_1_TQ[0]), .q(N31P_1_2P_1_STATES[1]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE), .gr(RESET_n));
xor2 N31P_1_2P_1_83P_1_I23_1_I8_1 (.o(N31P_1_2P_1_83P_1_I23_1_TQ[0]), .i0(N31P_1_2P_1_83P_1_T5), .i1(N31P_1_2P_1_STATES[5]));
fdce N31P_1_2P_1_83P_1_I23_1_I7_1 (.gr(XVDD), .d(N31P_1_2P_1_83P_1_I23_1_TQ[0]), .q(N31P_1_2P_1_STATES[5]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE));
xor2 N31P_1_2P_1_83P_1_I20_1_I8_1 (.o(N31P_1_2P_1_83P_1_I20_1_TQ[0]), .i0(N31P_1_2P_1_83P_1_T2), .i1(N31P_1_2P_1_STATES[2]));
fdce N31P_1_2P_1_83P_1_I20_1_I7_1 (.d(N31P_1_2P_1_83P_1_I20_1_TQ[0]), .q(N31P_1_2P_1_STATES[2]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE), .gr(RESET_n));
xor2 N31P_1_2P_1_83P_1_I18_1_I8_1 (.o(N31P_1_2P_1_83P_1_I18_1_TQ[0]), .i0(N31P_1_2P_1_83P_1_T3), .i1(N31P_1_2P_1_STATES[3]));
fdce N31P_1_2P_1_83P_1_I18_1_I7_1 (.d(N31P_1_2P_1_83P_1_I18_1_TQ[0]), .q(N31P_1_2P_1_STATES[3]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE), .gr(RESET_n));
xor2 N31P_1_2P_1_83P_1_I15_1_I8_1 (.o(N31P_1_2P_1_83P_1_I15_1_TQ[0]), .i0(N31P_1_2P_1_83P_1_T7), .i1(N31P_1_2P_1_STATES[7]));
fdce N31P_1_2P_1_83P_1_I15_1_I7_1 (.gr(XVDD), .d(N31P_1_2P_1_83P_1_I15_1_TQ[0]), .q(N31P_1_2P_1_STATES[7]), .c(CLK), .ce(N31P_1_2P_1_STAGE_ENABLE), .clr(N31P_1_2P_1_STAGE_DONE));
and3 N31P_1_2P_1_83P_1_I33_1 (.i2(N31P_1_2P_1_83P_1_T4), .o(N31P_1_2P_1_83P_1_T6), .i0(N31P_1_2P_1_STATES[5]), .i1(N31P_1_2P_1_STATES[4]));
and3 N31P_1_2P_1_83P_1_I32_1 (.i2(N31P_1_2P_1_STATES[0]), .o(N31P_1_2P_1_83P_1_T3), .i0(N31P_1_2P_1_STATES[2]), .i1(N31P_1_2P_1_STATES[1]));
and5 N31P_1_2P_1_83P_1_I25_1 (.i4(N31P_1_2P_1_83P_1_T4), .i2(N31P_1_2P_1_STATES[5]), .i3(N31P_1_2P_1_STATES[4]), .o(N31P_1_2P_1_83P_1_TC), .i0(N31P_1_2P_1_STATES[7]), .i1(N31P_1_2P_1_STATES[6]));
and4 N31P_1_2P_1_83P_1_I24_1 (.i2(N31P_1_2P_1_STATES[4]), .i3(N31P_1_2P_1_83P_1_T4), .o(N31P_1_2P_1_83P_1_T7), .i0(N31P_1_2P_1_STATES[6]), .i1(N31P_1_2P_1_STATES[5]));
and4 N31P_1_2P_1_83P_1_I16_1 (.i2(N31P_1_2P_1_STATES[1]), .i3(N31P_1_2P_1_STATES[0]), .o(N31P_1_2P_1_83P_1_T4), .i0(N31P_1_2P_1_STATES[3]), .i1(N31P_1_2P_1_STATES[2]));
and2 N31P_1_2P_1_83P_1_I29_1 (.o(N31P_1_2P_1_83P_1_T2), .i0(N31P_1_2P_1_STATES[1]), .i1(N31P_1_2P_1_STATES[0]));
and2 N31P_1_2P_1_83P_1_I22_1 (.o(N31P_1_2P_1_83P_1_CEO), .i0(N31P_1_2P_1_STAGE_ENABLE), .i1(N31P_1_2P_1_83P_1_TC));
and2 N31P_1_2P_1_83P_1_I21_1 (.o(N31P_1_2P_1_83P_1_T5), .i0(N31P_1_2P_1_STATES[4]), .i1(N31P_1_2P_1_83P_1_T4));
fdce N31P_1_2P_1_69P_1_I8_1 (.d(XVDD), .q(N31P_1_2P_1_STAGE_ENABLE), .c(N31P_1_2P_1_A), .ce(XVDD), .clr(N31P_1_CMOS_END), .gr(RESET_n));
inv N31P_1_2P_1_77P_1_21P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_21P_I), .o(N31P_1_2P_1_77P_1_UN_1_INV_20P_I));
inv N31P_1_2P_1_77P_1_22P_1 (.i(N31P_1_2P_1_CMOS_OP), .o(N31P_1_2P_1_77P_1_UN_1_INV_21P_I));
inv N31P_1_2P_1_77P_1_20P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_20P_I), .o(N31P_1_2P_1_77P_1_UN_1_INV_14P_I));
inv N31P_1_2P_1_77P_1_19P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_18P_O), .o(N31P_1_2P_1_77P_1_UN_1_INV_13P_I));
inv N31P_1_2P_1_77P_1_18P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_17P_O), .o(N31P_1_2P_1_77P_1_UN_1_INV_18P_O));
inv N31P_1_2P_1_77P_1_17P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_16P_O), .o(N31P_1_2P_1_77P_1_UN_1_INV_17P_O));
inv N31P_1_2P_1_77P_1_16P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_15P_O), .o(N31P_1_2P_1_77P_1_UN_1_INV_16P_O));
inv N31P_1_2P_1_77P_1_15P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_14P_O), .o(N31P_1_2P_1_77P_1_UN_1_INV_15P_O));
inv N31P_1_2P_1_77P_1_14P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_14P_I), .o(N31P_1_2P_1_77P_1_UN_1_INV_14P_O));
inv N31P_1_2P_1_77P_1_13P_1 (.i(N31P_1_2P_1_77P_1_UN_1_INV_13P_I), .o(N31P_1_2P_1_CMOS_OP_DELAY));
inv N31P_1_2P_1_46P_1_21P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_21P_I), .o(N31P_1_2P_1_46P_1_UN_1_INV_20P_I));
inv N31P_1_2P_1_46P_1_22P_1 (.i(N31P_1_2P_1_STAGE_ENABLE), .o(N31P_1_2P_1_46P_1_UN_1_INV_21P_I));
inv N31P_1_2P_1_46P_1_20P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_20P_I), .o(N31P_1_2P_1_46P_1_UN_1_INV_14P_I));
inv N31P_1_2P_1_46P_1_19P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_18P_O), .o(N31P_1_2P_1_46P_1_UN_1_INV_13P_I));
inv N31P_1_2P_1_46P_1_18P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_17P_O), .o(N31P_1_2P_1_46P_1_UN_1_INV_18P_O));
inv N31P_1_2P_1_46P_1_17P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_16P_O), .o(N31P_1_2P_1_46P_1_UN_1_INV_17P_O));
inv N31P_1_2P_1_46P_1_16P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_15P_O), .o(N31P_1_2P_1_46P_1_UN_1_INV_16P_O));
inv N31P_1_2P_1_46P_1_15P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_14P_O), .o(N31P_1_2P_1_46P_1_UN_1_INV_15P_O));
inv N31P_1_2P_1_46P_1_14P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_14P_I), .o(N31P_1_2P_1_46P_1_UN_1_INV_14P_O));
inv N31P_1_2P_1_46P_1_13P_1 (.i(N31P_1_2P_1_46P_1_UN_1_INV_13P_I), .o(ACCESS_CMOS));
and5 N31P_1_2P_1_88P_1 (.i4(N31P_1_2P_1_STATES[0]), .i2(N31P_1_2P_1_STATES[2]), .i3(N31P_1_2P_1_STATES[1]), .o(N31P_1_CMOS_END), .i0(N31P_1_2P_1_UN_1_D3_8E_51P_E), .i1(N31P_1_2P_1_STATES[3]));
and2b2 N31P_1_2P_1_54P_1 (.o(N31P_1_2P_1_UN_1_D3_8E_52P_E), .i1(N31P_1_2P_1_CMOS_OP), .i0(N31P_1_2P_1_STATES[4]));
xor2 N31P_1_2P_1_42P_1 (.o(N31P_1_2P_1_UN_1_NAND2_41P_I0), .i0(N31P_1_2P_1_STATES[1]), .i1(N31P_1_2P_1_STATES[0]));
nand2 N31P_1_2P_1_41P_1 (.o(RD_STROBE_n), .i0(N31P_1_2P_1_UN_1_NAND2_41P_I0), .i1(N31P_1_2P_1_CMOS_DIG_ACCESS));
or2 N31P_1_2P_1_56P_1 (.o(N31P_1_2P_1_A), .i0(CADD_ENABLE), .i1(N31P_1_2P_1_REAL_DATA));
or2 N31P_1_2P_1_53P_1 (.o(N31P_1_2P_1_UN_1_D3_8E_51P_E), .i0(N31P_1_2P_1_CMOS_OP), .i1(N31P_1_2P_1_STATES[4]));
or2 N31P_1_2P_1_16P_1 (.o(N31P_1_2P_1_UN_1_OR2_16P_O), .i0(LATCH[2]), .i1(N31P_1_2P_1_STROBE[2]));
or2 N31P_1_2P_1_15P_1 (.o(N31P_1_2P_1_UN_1_OR2_15P_O), .i0(LATCH[3]), .i1(N31P_1_2P_1_STROBE[3]));
or2 N31P_1_2P_1_14P_1 (.o(N31P_1_2P_1_UN_1_OR2_14P_O), .i0(LATCH[4]), .i1(N31P_1_2P_1_STROBE[4]));
or2 N31P_1_2P_1_13P_1 (.o(N31P_1_2P_1_UN_1_OR2_13P_O), .i0(LATCH[1]), .i1(N31P_1_2P_1_STROBE[1]));
or4 N31P_1_2P_1_29P_1 (.i2(N31P_1_2P_1_UN_1_OR2_16P_O), .i3(N31P_1_2P_1_UN_1_OR2_13P_O), .o(N31P_1_2P_1_CMOS_DIG_ACCESS), .i0(N31P_1_2P_1_UN_1_OR2_14P_O), .i1(N31P_1_2P_1_UN_1_OR2_15P_O));
and2b1 N31P_1_2P_1_76P_1 (.o(N31P_1_2P_1_STAGE_DONE), .i0(ADC_BUSY), .i1(N31P_1_CMOS_END));
and2b1 N31P_1_2P_1_72P_1 (.o(N31P_1_DATA_READY), .i0(N31P_1_2P_1_CMOS_OP_DELAY), .i1(N31P_1_2P_1_STAGE_DONE));
and2 N31P_1_2P_1_79P_1 (.o(N31P_1_2P_1_REAL_DATA), .i0(N31P_1_ALL_DATA_PROCESSED), .i1(DATA_AVAILABLE));
inv N31P_1_2P_1_82P_1 (.i(CADD_ENABLE), .o(N31P_1_2P_1_UN_1_INV_81P_I));
inv N31P_1_2P_1_81P_1 (.i(N31P_1_2P_1_UN_1_INV_81P_I), .o(N31P_1_2P_1_CMOS_OP));
and3b1 N31P_1_9P_1 (.i2(LATCH_TAG), .o(GET_DATA), .i0(CREG_REQ), .i1(N31P_1_ALL_DATA_PROCESSED));
inv N31P_1_46P_1 (.i(N31P_1_UN_1_FDC_42P_Q), .o(CMOSR_DTACK_n));
inv N31P_1_45P_1 (.i(CADD_ENABLE), .o(N31P_1_UN_1_INV_44P_I));
inv N31P_1_44P_1 (.i(N31P_1_UN_1_INV_44P_I), .o(CREG_SEL));
bufg N70P_1 (.i(SQCLK), .o(CLK));
bufg N69P_1 (.i(UN_1_BUFG_69P_I), .o(CLKD2));
and2 N82P_1_3 (.o(UN_1_AND2_82P_O[2]), .i0(UN_1_AND2_82P_I0[2]), .i1(UN_1_AND2_82P_I0[2]));
and2 N82P_1_2 (.i1(UN_1_AND2_82P_I0[1]), .i0(UN_1_AND2_82P_I0[1]), .o(UN_1_AND2_82P_O[1]));
and2 N82P_1_1 (.i1(UN_1_AND2_82P_I0[0]), .i0(UN_1_AND2_82P_I0[0]), .o(UN_1_AND2_82P_O[0]));
and2 N54P_1 (.o(UN_1_AND2_54P_O), .i0(UN_1_AND2_54P_I0), .i1(UN_1_AND2_54P_I0));
ibuf N83P_1_3 (.i(SPAREIN[2]), .o(UN_1_AND2_82P_I0[2]));
ibuf N83P_1_2 (.o(UN_1_AND2_82P_I0[1]), .i(SPAREIN[1]));
ibuf N83P_1_1 (.o(UN_1_AND2_82P_I0[0]), .i(SPAREIN[0]));
ibuf N45P_1_3 (.i(SQXREG_SEL[2]), .o(REG_SEL[2]));
ibuf N45P_1_2 (.o(REG_SEL[1]), .i(SQXREG_SEL[1]));
ibuf N45P_1_1 (.o(REG_SEL[0]), .i(SQXREG_SEL[0]));
ibuf N73P_1 (.i(SQADC_BUSY_n), .o(UN_1_IBUF_73P_O));
ibuf N72P_1 (.i(SQMEMORY_ACK_n), .o(MEMORY_ACK_n));
ibuf N53P_1 (.i(SDIN), .o(UN_1_AND2_54P_I0));
ibuf N49P_1 (.i(SQXREG_RD_n), .o(REG_RD_n));
ibuf N48P_1 (.i(SQXREG_WR_n), .o(REG_WR_n));
inv N57P_1 (.i(GET_DATA), .o(UN_1_INV_57P_O));
inv N34P_1 (.i(UN_1_IBUF_73P_O), .o(ADC_BUSY));
inv N33P_1 (.i(CONVERT_START), .o(UN_1_INV_33P_O));
obuf N76P_1_5 (.i(TAG[4]), .o(SQTAG[4]));
obuf N76P_1_4 (.o(SQTAG[3]), .i(TAG[3]));
obuf N76P_1_3 (.o(SQTAG[2]), .i(TAG[2]));
obuf N76P_1_2 (.o(SQTAG[1]), .i(TAG[1]));
obuf N76P_1_1 (.o(SQTAG[0]), .i(TAG[0]));
obuf N12P_1_4 (.i(LATCH[4]), .o(SQLATCH[4]));
obuf N12P_1_3 (.o(SQLATCH[3]), .i(LATCH[3]));
obuf N12P_1_2 (.o(SQLATCH[2]), .i(LATCH[2]));
obuf N12P_1_1 (.o(SQLATCH[1]), .i(LATCH[1]));
obuf N80P_1_3 (.i(UN_1_AND2_82P_O[2]), .o(SPAREOUT[2]));
obuf N80P_1_2 (.o(SPAREOUT[1]), .i(UN_1_AND2_82P_O[1]));
obuf N80P_1_1 (.o(SPAREOUT[0]), .i(UN_1_AND2_82P_O[0]));
obuf N10P_1_3 (.i(ENW_[3]), .o(SQENW_[3]));
obuf N10P_1_2 (.o(SQENW_[2]), .i(ENW_[2]));
obuf N10P_1_1 (.o(SQENW_[1]), .i(ENW_[1]));
obuf N78P_1 (.i(XVDD), .o(ADC_DONE));
obuf N75P_1 (.i(CMOSR_DTACK_n), .o(SQCHOLD_n));
obuf N63P_1 (.i(CREG_SEL), .o(SQCREG_SEL));
obuf N61P_1 (.i(ACCESS_CMOS), .o(SQCHIP_SEL_EN));
obuf N59P_1 (.i(UN_1_INV_57P_O), .o(SQFECBUSY));
obuf N56P_1 (.i(UN_1_AND2_54P_O), .o(SDOUT));
obuf N51P_1 (.i(XVDD), .o(M2));
obuf N29P_1 (.i(DAV32OR), .o(SQDAV32OR));
obuf N14P_1 (.i(UN_1_INV_33P_O), .o(SQCONVERT_START_n));
obuf N13P_1 (.i(RD_STROBE_n), .o(SQRD_STROBE_n));
obuf N11P_1 (.i(MEMORY_REQUEST_n), .o(SQMEMORY_REQUEST_n));
obuf N9P_1 (.i(CADD_ENABLE), .o(SQCADD_ENABLE));
endmodule
`uselib

module seq96new_globals();

wire GR;
endmodule

