/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from xcountsynct.xcd on Fri Sep 20 01:21:40 1996 */
/* PART 3190PQ160-3 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module xcountsynct
(X50MHZ, X10MHZ, XTRIGCOMB, XTC_24_n, XTC_16_n, XSYNCLR24, xsynclr, XSYNC, xspecial_raw, XRESYNC, XLOCKOUT_n, XLOAD_SYNC50_n, XLOAD_SYNC10_n, XLOAD_EN50_n, XLOAD_EN10_n, XLOAD_ENGT_n, XGTRIG, XGTLOAD24_n, XGTLOAD16_n, XGTCLK24, XGTCLK16, XGCLK, XFF_LA, XERR, XEF_LA, XCLK_SYNC10, XASYNC_EN, SPARES, SDOUT, SDIN, M2, RESET_n, DUMMY_OUT, RDATA_n, RTRIG, PROGRAM_n, CCLK, PWRDWN_n);
   input X50MHZ;
   input X10MHZ;
   input [8:0] XTRIGCOMB;
   input XTC_24_n;
   input XTC_16_n;
   output XSYNCLR24;
   output xsynclr;
   input XSYNC;
   output xspecial_raw;
   input XRESYNC;
   input XLOCKOUT_n;
   output XLOAD_SYNC50_n;
   output XLOAD_SYNC10_n;
   input XLOAD_EN50_n;
   input XLOAD_EN10_n;
   input XLOAD_ENGT_n;
   input XGTRIG;
   output XGTLOAD24_n;
   output XGTLOAD16_n;
   output XGTCLK24;
   output XGTCLK16;
   output XGCLK;
   input [23:0] XFF_LA;
   output [6:0] XERR;
   input [23:0] XEF_LA;
   output XCLK_SYNC10;
   input XASYNC_EN;
   input [9:0] SPARES;
   output SDOUT;
   input SDIN;
   output M2;
   input RESET_n;
   output DUMMY_OUT;
   output RDATA_n;
   input RTRIG;
   input PROGRAM_n;
   input CCLK;
   input PWRDWN_n;
wire [0:0] N60P_1_10P_1_I35;
wire [0:0] N48P_1_27P_1_38P_1_I47;
wire [0:0] N48P_1_27P_1_32P_1_I47;
wire [0:0] N48P_1_27P_1_31P_1_I47;
wire [0:0] N48P_1_27P_1_30P_1_I47;
wire [0:0] N48P_1_27P_1_29P_1_I47;
wire [0:0] N48P_1_27P_1_28P_1_I47;
wire [0:0] N48P_1_26P_1_38P_1_I47;
wire [0:0] N48P_1_26P_1_32P_1_I47;
wire [0:0] N48P_1_26P_1_31P_1_I47;
wire [0:0] N48P_1_26P_1_30P_1_I47;
wire [0:0] N48P_1_26P_1_29P_1_I47;
wire [0:0] N48P_1_26P_1_28P_1_I47;
wire [4:0] UN_1_IBUF_67P_O;
wire [8:0] TRIGCOMB;
wire [23:0] FF_LA;
wire [6:0] ERR;
wire [23:0] EF_LA;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/neubauer/xilinx/xcountsynct/verilog_lib/xcountsynct.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

and4 N60P_1_10P_1_I11_1 (.i0(TRIGCOMB[2]), .i1(TRIGCOMB[3]), .i2(TRIGCOMB[5]), .i3(N60P_1_10P_1_I35[0]), .o(UN_1_OBUF_64P_I));
and3 N60P_1_10P_1_I8_1 (.i0(TRIGCOMB[6]), .i1(TRIGCOMB[7]), .i2(TRIGCOMB[8]), .o(N60P_1_10P_1_I35[0]));
and3 N60P_1_8P_1 (.i0(TRIGCOMB[0]), .i1(N60P_1_UN_1_AND3_8P_I1), .i2(TRIGCOMB[4]), .o(SPECIAL_RAW));
inv N60P_1_2P_1 (.i(TRIGCOMB[1]), .o(N60P_1_UN_1_AND3_8P_I1));
fdce N5P_1_3P_1_I8_1 (.q(N5P_1_UN_1_FDC_3P_Q), .d(XVDD), .c(N5P_1_UN_1_AND2_6P_O), .ce(XVDD), .clr(N5P_1_UN_1_AND2_5P_O), .gr(RESET_n));
fdce N5P_1_4P_1_I8_1 (.q(N5P_1_UN_1_AND2_6P_I0), .d(XVDD), .c(GTRIG_ACLK), .ce(XVDD), .clr(N5P_1_UN_1_AND2_5P_I0), .gr(RESET_n));
inv N5P_1_8P_1 (.i(gclk), .o(N5P_1_UN_1_INV_8P_O));
inv N5P_1_9P_1 (.i(N5P_1_UN_1_INV_8P_O), .o(N5P_1_UN_1_AND2_5P_I0));
inv N5P_1_13P_1 (.i(N5P_1_UN_1_INV_12P_O), .o(gclk));
inv N5P_1_12P_1 (.i(N5P_1_UN_1_INV_11P_O), .o(N5P_1_UN_1_INV_12P_O));
inv N5P_1_11P_1 (.i(N5P_1_UN_1_INV_10P_O), .o(N5P_1_UN_1_INV_11P_O));
inv N5P_1_10P_1 (.i(N5P_1_UN_1_FDC_3P_Q), .o(N5P_1_UN_1_INV_10P_O));
and2 N5P_1_5P_1 (.i0(N5P_1_UN_1_AND2_5P_I0), .i1(N10MHZ), .o(N5P_1_UN_1_AND2_5P_O));
and2 N5P_1_6P_1 (.i0(N5P_1_UN_1_AND2_6P_I0), .i1(N10MHZ), .o(N5P_1_UN_1_AND2_6P_O));
fdce N4P_1_45P_1_I8_1 (.q(N4P_1_UN_1_AND2_44P_I1), .d(XVDD), .c(SYNCLR), .ce(XVDD), .clr(N4P_1_CLR16), .gr(RESET_n));
fdce N4P_1_41P_1_I8_1 (.q(N4P_1_UN_1_AND2_42P_I1), .d(XVDD), .c(SYNCLR24), .ce(XVDD), .clr(N4P_1_CLR24), .gr(RESET_n));
or2 N4P_1_36P_1 (.i0(N4P_1_CLR24), .i1(GTRIG), .o(GTCLK24));
or2 N4P_1_18P_1 (.i0(GTRIG), .i1(N4P_1_CLR16), .o(GTCLK16));
inv N4P_1_43P_1 (.i(N4P_1_UN_1_AND2_42P_I1), .o(GTLOAD24_n));
inv N4P_1_39P_1 (.i(N4P_1_UN_1_AND2_44P_I1), .o(GTLOAD16_n));
and2 N4P_1_44P_1 (.i0(LOCKOUT_n), .i1(N4P_1_UN_1_AND2_44P_I1), .o(N4P_1_CLR16));
and2 N4P_1_42P_1 (.i0(LOCKOUT_n), .i1(N4P_1_UN_1_AND2_42P_I1), .o(N4P_1_CLR24));
fdce N48P_1_13P_1_I8_1 (.q(ERR[0]), .d(XVDD), .c(SYNCLR), .ce(XVDD), .clr(LOCKOUT_n), .gr(RESET_n));
fdce N48P_1_12P_1_I8_1 (.q(N48P_1_UN_1_FDC_12P_Q), .d(XVDD), .c(N48P_1_UN_1_FDC_12P_C), .ce(XVDD), .clr(LOCKOUT_n), .gr(RESET_n));
fdce N48P_1_11P_1_I8_1 (.q(ERR[2]), .d(XVDD), .c(SYNCLR24), .ce(XVDD), .clr(LOCKOUT_n), .gr(RESET_n));
fdce N48P_1_10P_1_I8_1 (.q(N48P_1_UN_1_FDC_10P_Q), .d(XVDD), .c(N48P_1_UN_1_FDC_10P_C), .ce(XVDD), .clr(LOCKOUT_n), .gr(RESET_n));
nand5 N48P_1_27P_1_38P_1_I10_1 (.i0(FF_LA[16]), .i1(FF_LA[17]), .i2(FF_LA[18]), .i3(FF_LA[19]), .i4(N48P_1_27P_1_38P_1_I47[0]), .o(N48P_1_27P_1_UN_1_NAND8_38P_O));
and4 N48P_1_27P_1_38P_1_I12_1 (.i0(FF_LA[20]), .i1(FF_LA[21]), .i2(FF_LA[22]), .i3(FF_LA[23]), .o(N48P_1_27P_1_38P_1_I47[0]));
nand5 N48P_1_27P_1_32P_1_I10_1 (.i0(FF_LA[8]), .i1(FF_LA[9]), .i2(FF_LA[10]), .i3(FF_LA[11]), .i4(N48P_1_27P_1_32P_1_I47[0]), .o(N48P_1_27P_1_UN_1_NAND8_32P_O));
and4 N48P_1_27P_1_32P_1_I12_1 (.i0(FF_LA[12]), .i1(FF_LA[13]), .i2(FF_LA[14]), .i3(FF_LA[15]), .o(N48P_1_27P_1_32P_1_I47[0]));
nand5 N48P_1_27P_1_31P_1_I10_1 (.i0(FF_LA[0]), .i1(FF_LA[1]), .i2(FF_LA[2]), .i3(FF_LA[3]), .i4(N48P_1_27P_1_31P_1_I47[0]), .o(N48P_1_27P_1_UN_1_NAND8_31P_O));
and4 N48P_1_27P_1_31P_1_I12_1 (.i0(FF_LA[4]), .i1(FF_LA[5]), .i2(FF_LA[6]), .i3(FF_LA[7]), .o(N48P_1_27P_1_31P_1_I47[0]));
or5 N48P_1_27P_1_30P_1_I10_1 (.i0(FF_LA[16]), .i1(FF_LA[17]), .i2(FF_LA[18]), .i3(FF_LA[19]), .i4(N48P_1_27P_1_30P_1_I47[0]), .o(N48P_1_27P_1_UN_1_OR3_27P_I2));
or4 N48P_1_27P_1_30P_1_I13_1 (.i0(FF_LA[20]), .i1(FF_LA[21]), .i2(FF_LA[22]), .i3(FF_LA[23]), .o(N48P_1_27P_1_30P_1_I47[0]));
or5 N48P_1_27P_1_29P_1_I10_1 (.i0(FF_LA[8]), .i1(FF_LA[9]), .i2(FF_LA[10]), .i3(FF_LA[11]), .i4(N48P_1_27P_1_29P_1_I47[0]), .o(N48P_1_27P_1_UN_1_OR3_27P_I1));
or4 N48P_1_27P_1_29P_1_I13_1 (.i0(FF_LA[12]), .i1(FF_LA[13]), .i2(FF_LA[14]), .i3(FF_LA[15]), .o(N48P_1_27P_1_29P_1_I47[0]));
or5 N48P_1_27P_1_28P_1_I10_1 (.i0(FF_LA[0]), .i1(FF_LA[1]), .i2(FF_LA[2]), .i3(FF_LA[3]), .i4(N48P_1_27P_1_28P_1_I47[0]), .o(N48P_1_27P_1_UN_1_OR3_27P_I0));
or4 N48P_1_27P_1_28P_1_I13_1 (.i0(FF_LA[4]), .i1(FF_LA[5]), .i2(FF_LA[6]), .i3(FF_LA[7]), .o(N48P_1_27P_1_28P_1_I47[0]));
inv N48P_1_27P_1_41P_1 (.i(N48P_1_27P_1_ALL_LOW_n), .o(ERR[6]));
and2 N48P_1_27P_1_24P_1 (.i0(N48P_1_27P_1_ALL_HIGH_n), .i1(N48P_1_27P_1_ALL_LOW_n), .o(ERR[5]));
or3 N48P_1_27P_1_27P_1 (.i0(N48P_1_27P_1_UN_1_OR3_27P_I0), .i1(N48P_1_27P_1_UN_1_OR3_27P_I1), .i2(N48P_1_27P_1_UN_1_OR3_27P_I2), .o(N48P_1_27P_1_ALL_LOW_n));
or3 N48P_1_27P_1_26P_1 (.i0(N48P_1_27P_1_UN_1_NAND8_31P_O), .i1(N48P_1_27P_1_UN_1_NAND8_32P_O), .i2(N48P_1_27P_1_UN_1_NAND8_38P_O), .o(N48P_1_27P_1_ALL_HIGH_n));
nand5 N48P_1_26P_1_38P_1_I10_1 (.i0(EF_LA[16]), .i1(EF_LA[17]), .i2(EF_LA[18]), .i3(EF_LA[19]), .i4(N48P_1_26P_1_38P_1_I47[0]), .o(N48P_1_26P_1_UN_1_NAND8_38P_O));
and4 N48P_1_26P_1_38P_1_I12_1 (.i0(EF_LA[20]), .i1(EF_LA[21]), .i2(EF_LA[22]), .i3(EF_LA[23]), .o(N48P_1_26P_1_38P_1_I47[0]));
nand5 N48P_1_26P_1_32P_1_I10_1 (.i0(EF_LA[8]), .i1(EF_LA[9]), .i2(EF_LA[10]), .i3(EF_LA[11]), .i4(N48P_1_26P_1_32P_1_I47[0]), .o(N48P_1_26P_1_UN_1_NAND8_32P_O));
and4 N48P_1_26P_1_32P_1_I12_1 (.i0(EF_LA[12]), .i1(EF_LA[13]), .i2(EF_LA[14]), .i3(EF_LA[15]), .o(N48P_1_26P_1_32P_1_I47[0]));
nand5 N48P_1_26P_1_31P_1_I10_1 (.i0(EF_LA[0]), .i1(EF_LA[1]), .i2(EF_LA[2]), .i3(EF_LA[3]), .i4(N48P_1_26P_1_31P_1_I47[0]), .o(N48P_1_26P_1_UN_1_NAND8_31P_O));
and4 N48P_1_26P_1_31P_1_I12_1 (.i0(EF_LA[4]), .i1(EF_LA[5]), .i2(EF_LA[6]), .i3(EF_LA[7]), .o(N48P_1_26P_1_31P_1_I47[0]));
or5 N48P_1_26P_1_30P_1_I10_1 (.i0(EF_LA[16]), .i1(EF_LA[17]), .i2(EF_LA[18]), .i3(EF_LA[19]), .i4(N48P_1_26P_1_30P_1_I47[0]), .o(N48P_1_26P_1_UN_1_OR3_27P_I2));
or4 N48P_1_26P_1_30P_1_I13_1 (.i0(EF_LA[20]), .i1(EF_LA[21]), .i2(EF_LA[22]), .i3(EF_LA[23]), .o(N48P_1_26P_1_30P_1_I47[0]));
or5 N48P_1_26P_1_29P_1_I10_1 (.i0(EF_LA[8]), .i1(EF_LA[9]), .i2(EF_LA[10]), .i3(EF_LA[11]), .i4(N48P_1_26P_1_29P_1_I47[0]), .o(N48P_1_26P_1_UN_1_OR3_27P_I1));
or4 N48P_1_26P_1_29P_1_I13_1 (.i0(EF_LA[12]), .i1(EF_LA[13]), .i2(EF_LA[14]), .i3(EF_LA[15]), .o(N48P_1_26P_1_29P_1_I47[0]));
or5 N48P_1_26P_1_28P_1_I10_1 (.i0(EF_LA[0]), .i1(EF_LA[1]), .i2(EF_LA[2]), .i3(EF_LA[3]), .i4(N48P_1_26P_1_28P_1_I47[0]), .o(N48P_1_26P_1_UN_1_OR3_27P_I0));
or4 N48P_1_26P_1_28P_1_I13_1 (.i0(EF_LA[4]), .i1(EF_LA[5]), .i2(EF_LA[6]), .i3(EF_LA[7]), .o(N48P_1_26P_1_28P_1_I47[0]));
inv N48P_1_26P_1_41P_1 (.i(N48P_1_26P_1_ALL_LOW_n), .o(N48P_1_26P_1_ALL_LOW));
and2 N48P_1_26P_1_24P_1 (.i0(N48P_1_26P_1_ALL_HIGH_n), .i1(N48P_1_26P_1_ALL_LOW_n), .o(ERR[4]));
or3 N48P_1_26P_1_27P_1 (.i0(N48P_1_26P_1_UN_1_OR3_27P_I0), .i1(N48P_1_26P_1_UN_1_OR3_27P_I1), .i2(N48P_1_26P_1_UN_1_OR3_27P_I2), .o(N48P_1_26P_1_ALL_LOW_n));
or3 N48P_1_26P_1_26P_1 (.i0(N48P_1_26P_1_UN_1_NAND8_31P_O), .i1(N48P_1_26P_1_UN_1_NAND8_32P_O), .i2(N48P_1_26P_1_UN_1_NAND8_38P_O), .o(N48P_1_26P_1_ALL_HIGH_n));
inv N48P_1_31P_1 (.i(TC_16_n), .o(N48P_1_UN_1_FDC_12P_C));
inv N48P_1_30P_1 (.i(TC_24_n), .o(N48P_1_UN_1_FDC_10P_C));
xor2 N48P_1_32P_1 (.i0(N48P_1_UN_1_FDC_10P_Q), .i1(ERR[2]), .o(ERR[3]));
xor2 N48P_1_33P_1 (.i0(N48P_1_UN_1_FDC_12P_Q), .i1(ERR[0]), .o(ERR[1]));
fdce N2P_1_8P_1_I6_1 (.q(N2P_1_UN_1_FDC_1_8P_Q), .d(XVDD), .c(N2P_1_8P_1_CB), .ce(XVDD), .clr(N2P_1_UN_1_FDC_1_8P_CLR), .gr(RESET_n));
inv N2P_1_8P_1_I7_1 (.i(LOAD_EN10_n), .o(N2P_1_8P_1_CB));
or2 N2P_1_11P_1 (.i0(N2P_1_UN_1_AND2_10P_O), .i1(SYNC), .o(CLK_SYNC10));
inv N2P_1_6P_1 (.i(SYNC), .o(N2P_1_UN_1_INV_6P_O));
inv N2P_1_7P_1 (.i(N2P_1_UN_1_INV_6P_O), .o(N2P_1_UN_1_FDC_1_8P_CLR));
inv N2P_1_9P_1 (.i(N2P_1_UN_1_FDC_1_8P_Q), .o(LOAD_SYNC10_n));
and2 N2P_1_10P_1 (.i0(LOAD_SYNC10_n), .i1(N10MHZ), .o(N2P_1_UN_1_AND2_10P_O));
fdce N1P_1_6P_1_I8_1 (.q(N1P_1_UN_1_FDC_6P_Q), .d(XVDD), .c(N1P_1_UN_1_AND2_5P_O), .ce(XVDD), .clr(N1P_1_UN_1_FDC_6P_CLR), .gr(RESET_n));
or2 N1P_1_4P_1 (.i0(N1P_1_UN_1_FDC_6P_Q), .i1(LOAD_EN50_n), .o(LOAD_SYNC50_n));
inv N1P_1_7P_1 (.i(N1P_1_UN_1_AND2_5P_I1), .o(N1P_1_UN_1_FDC_6P_CLR));
inv N1P_1_8P_1 (.i(LOAD_EN50_n), .o(N1P_1_UN_1_AND2_5P_I1));
and2 N1P_1_5P_1 (.i0(N50MHZ), .i1(N1P_1_UN_1_AND2_5P_I1), .o(N1P_1_UN_1_AND2_5P_O));
fdce N3P_1_83P_1_I6_1 (.q(N3P_1_SYNC24RS), .d(N3P_1_UN_1_FD_82P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_82P_1_I6_1 (.q(N3P_1_UN_1_FD_82P_Q), .d(N3P_1_UN_1_FD_81P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_81P_1_I6_1 (.q(N3P_1_UN_1_FD_81P_Q), .d(N3P_1_UN_1_FD_80P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_80P_1_I6_1 (.q(N3P_1_UN_1_FD_80P_Q), .d(N3P_1_UN_1_FD_79P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_79P_1_I6_1 (.q(N3P_1_UN_1_FD_79P_Q), .d(SYNCLR24), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_76P_1_I6_1 (.q(N3P_1_SYNC16RS), .d(N3P_1_UN_1_FD_75P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_75P_1_I6_1 (.q(N3P_1_UN_1_FD_75P_Q), .d(N3P_1_UN_1_FD_74P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_74P_1_I6_1 (.q(N3P_1_UN_1_FD_74P_Q), .d(N3P_1_UN_1_FD_73P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_73P_1_I6_1 (.q(N3P_1_UN_1_FD_73P_Q), .d(N3P_1_UN_1_FD_72P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_72P_1_I6_1 (.q(N3P_1_UN_1_FD_72P_Q), .d(SYNCLR), .c(N50MHZ_GCLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_63P_1_I6_1 (.q(N3P_1_PRESET), .d(XVDD), .c(GTRIG_ACLK), .ce(XVDD), .clr(XGND), .gr(RESET_n));
fdce N3P_1_86P_1_I8_1 (.q(N3P_1_UN_1_AND2_41P_I1), .d(XVDD), .c(N3P_1_UN_1_FDC_86P_C), .ce(XVDD), .clr(N3P_1_SYNC16RS), .gr(RESET_n));
fdce N3P_1_85P_1_I8_1 (.q(N3P_1_UN_1_AND2_64P_I0), .d(XVDD), .c(N3P_1_UN_1_INV_59P_O), .ce(XVDD), .clr(N3P_1_SYNC24RS), .gr(RESET_n));
fdce N3P_1_84P_1_I8_1 (.q(N3P_1_UN_1_FDC_84P_Q), .d(XVDD), .c(N3P_1_UN_1_INV_67P_O), .ce(XVDD), .clr(N3P_1_SYNC16RS), .gr(RESET_n));
fdce N3P_1_71P_1_I8_1 (.q(SYNCLR), .d(N3P_1_UN_1_FDC_70P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(N3P_1_SYNC16RS), .gr(RESET_n));
fdce N3P_1_70P_1_I8_1 (.q(N3P_1_UN_1_FDC_70P_Q), .d(N3P_1_SYNC16), .c(N50MHZ_GCLK), .ce(XVDD), .clr(N3P_1_SYNC16RS), .gr(RESET_n));
fdce N3P_1_78P_1_I8_1 (.q(SYNCLR24), .d(N3P_1_UN_1_FDC_77P_Q), .c(N50MHZ_GCLK), .ce(XVDD), .clr(N3P_1_SYNC24RS), .gr(RESET_n));
fdce N3P_1_77P_1_I8_1 (.q(N3P_1_UN_1_FDC_77P_Q), .d(N3P_1_SYNC24), .c(N50MHZ_GCLK), .ce(XVDD), .clr(N3P_1_SYNC24RS), .gr(RESET_n));
inv N3P_1_67P_1 (.i(LOAD_ENGT_n), .o(N3P_1_UN_1_INV_67P_O));
inv N3P_1_59P_1 (.i(TC_24_n), .o(N3P_1_UN_1_INV_59P_O));
inv N3P_1_58P_1 (.i(TC_16_n), .o(N3P_1_UN_1_FDC_86P_C));
and2 N3P_1_65P_1 (.i0(N3P_1_PRESET), .i1(N3P_1_UN_1_AND2_41P_I1), .o(N3P_1_UN_1_AND2_65P_O));
and2 N3P_1_64P_1 (.i0(N3P_1_UN_1_AND2_64P_I0), .i1(N3P_1_PRESET), .o(N3P_1_UN_1_AND2_64P_O));
and2 N3P_1_41P_1 (.i0(RESYNC), .i1(N3P_1_UN_1_AND2_41P_I1), .o(N3P_1_UN_1_AND2_41P_O));
and2 N3P_1_16P_1 (.i0(GTRIG), .i1(ASYNC_EN), .o(N3P_1_UN_1_AND2_16P_O));
or3 N3P_1_69P_1 (.i0(N3P_1_UN_1_AND2_65P_O), .i1(N3P_1_UN_1_AND2_16P_O), .i2(N3P_1_UN_1_FDC_84P_Q), .o(N3P_1_SYNC16));
or4 N3P_1_66P_1 (.i0(N3P_1_UN_1_AND2_41P_O), .i1(N3P_1_UN_1_AND2_16P_O), .i2(N3P_1_UN_1_FDC_84P_Q), .i3(N3P_1_UN_1_AND2_64P_O), .o(N3P_1_SYNC24));
gclk N66P_1 (.i(N50MHZ), .o(N50MHZ_GCLK));
aclk N65P_1 (.i(GTRIG), .o(GTRIG_ACLK));
ibuf N58P_1_9 (.i(XTRIGCOMB[8]), .o(TRIGCOMB[8]));
ibuf N58P_1_8 (.o(TRIGCOMB[7]), .i(XTRIGCOMB[7]));
ibuf N58P_1_7 (.o(TRIGCOMB[6]), .i(XTRIGCOMB[6]));
ibuf N58P_1_6 (.o(TRIGCOMB[5]), .i(XTRIGCOMB[5]));
ibuf N58P_1_5 (.o(TRIGCOMB[4]), .i(XTRIGCOMB[4]));
ibuf N58P_1_4 (.o(TRIGCOMB[3]), .i(XTRIGCOMB[3]));
ibuf N58P_1_3 (.o(TRIGCOMB[2]), .i(XTRIGCOMB[2]));
ibuf N58P_1_2 (.o(TRIGCOMB[1]), .i(XTRIGCOMB[1]));
ibuf N58P_1_1 (.o(TRIGCOMB[0]), .i(XTRIGCOMB[0]));
ibuf N67P_1_5 (.i(SPARES[9]), .o(UN_1_IBUF_67P_O[4]));
ibuf N67P_1_4 (.o(UN_1_IBUF_67P_O[3]), .i(SPARES[8]));
ibuf N67P_1_3 (.o(UN_1_IBUF_67P_O[2]), .i(SPARES[7]));
ibuf N67P_1_2 (.o(UN_1_IBUF_67P_O[1]), .i(SPARES[6]));
ibuf N67P_1_1 (.o(UN_1_IBUF_67P_O[0]), .i(SPARES[5]));
ibuf N68P_1 (.i(SDIN), .o(UN_1_IBUF_68P_O));
ibuf N56P_1 (.i(XLOCKOUT_n), .o(LOCKOUT_n));
ibuf N32P_1 (.i(XLOAD_EN10_n), .o(LOAD_EN10_n));
ibuf N31P_1 (.i(XSYNC), .o(SYNC));
ibuf N30P_1 (.i(XLOAD_EN50_n), .o(LOAD_EN50_n));
ibuf N29P_1 (.i(XLOAD_ENGT_n), .o(LOAD_ENGT_n));
ibuf N28P_1 (.i(X50MHZ), .o(N50MHZ));
ibuf N27P_1 (.i(XGTRIG), .o(GTRIG));
ibuf N26P_1 (.i(XTC_16_n), .o(TC_16_n));
ibuf N25P_1 (.i(XTC_24_n), .o(TC_24_n));
ibuf N24P_1 (.i(XRESYNC), .o(RESYNC));
ibuf N23P_1 (.i(XASYNC_EN), .o(ASYNC_EN));
ibuf N33P_1 (.i(X10MHZ), .o(N10MHZ));
ibuf N53P_1_24 (.i(XEF_LA[23]), .o(EF_LA[23]));
ibuf N53P_1_23 (.o(EF_LA[22]), .i(XEF_LA[22]));
ibuf N53P_1_22 (.o(EF_LA[21]), .i(XEF_LA[21]));
ibuf N53P_1_21 (.o(EF_LA[20]), .i(XEF_LA[20]));
ibuf N53P_1_20 (.o(EF_LA[19]), .i(XEF_LA[19]));
ibuf N53P_1_19 (.o(EF_LA[18]), .i(XEF_LA[18]));
ibuf N53P_1_18 (.o(EF_LA[17]), .i(XEF_LA[17]));
ibuf N53P_1_17 (.o(EF_LA[16]), .i(XEF_LA[16]));
ibuf N53P_1_16 (.o(EF_LA[15]), .i(XEF_LA[15]));
ibuf N53P_1_15 (.o(EF_LA[14]), .i(XEF_LA[14]));
ibuf N53P_1_14 (.o(EF_LA[13]), .i(XEF_LA[13]));
ibuf N53P_1_13 (.o(EF_LA[12]), .i(XEF_LA[12]));
ibuf N53P_1_12 (.o(EF_LA[11]), .i(XEF_LA[11]));
ibuf N53P_1_11 (.o(EF_LA[10]), .i(XEF_LA[10]));
ibuf N53P_1_10 (.o(EF_LA[9]), .i(XEF_LA[9]));
ibuf N53P_1_9 (.o(EF_LA[8]), .i(XEF_LA[8]));
ibuf N53P_1_8 (.o(EF_LA[7]), .i(XEF_LA[7]));
ibuf N53P_1_7 (.o(EF_LA[6]), .i(XEF_LA[6]));
ibuf N53P_1_6 (.o(EF_LA[5]), .i(XEF_LA[5]));
ibuf N53P_1_5 (.o(EF_LA[4]), .i(XEF_LA[4]));
ibuf N53P_1_4 (.o(EF_LA[3]), .i(XEF_LA[3]));
ibuf N53P_1_3 (.o(EF_LA[2]), .i(XEF_LA[2]));
ibuf N53P_1_2 (.o(EF_LA[1]), .i(XEF_LA[1]));
ibuf N53P_1_1 (.o(EF_LA[0]), .i(XEF_LA[0]));
ibuf N51P_1_24 (.i(XFF_LA[23]), .o(FF_LA[23]));
ibuf N51P_1_23 (.o(FF_LA[22]), .i(XFF_LA[22]));
ibuf N51P_1_22 (.o(FF_LA[21]), .i(XFF_LA[21]));
ibuf N51P_1_21 (.o(FF_LA[20]), .i(XFF_LA[20]));
ibuf N51P_1_20 (.o(FF_LA[19]), .i(XFF_LA[19]));
ibuf N51P_1_19 (.o(FF_LA[18]), .i(XFF_LA[18]));
ibuf N51P_1_18 (.o(FF_LA[17]), .i(XFF_LA[17]));
ibuf N51P_1_17 (.o(FF_LA[16]), .i(XFF_LA[16]));
ibuf N51P_1_16 (.o(FF_LA[15]), .i(XFF_LA[15]));
ibuf N51P_1_15 (.o(FF_LA[14]), .i(XFF_LA[14]));
ibuf N51P_1_14 (.o(FF_LA[13]), .i(XFF_LA[13]));
ibuf N51P_1_13 (.o(FF_LA[12]), .i(XFF_LA[12]));
ibuf N51P_1_12 (.o(FF_LA[11]), .i(XFF_LA[11]));
ibuf N51P_1_11 (.o(FF_LA[10]), .i(XFF_LA[10]));
ibuf N51P_1_10 (.o(FF_LA[9]), .i(XFF_LA[9]));
ibuf N51P_1_9 (.o(FF_LA[8]), .i(XFF_LA[8]));
ibuf N51P_1_8 (.o(FF_LA[7]), .i(XFF_LA[7]));
ibuf N51P_1_7 (.o(FF_LA[6]), .i(XFF_LA[6]));
ibuf N51P_1_6 (.o(FF_LA[5]), .i(XFF_LA[5]));
ibuf N51P_1_5 (.o(FF_LA[4]), .i(XFF_LA[4]));
ibuf N51P_1_4 (.o(FF_LA[3]), .i(XFF_LA[3]));
ibuf N51P_1_3 (.o(FF_LA[2]), .i(XFF_LA[2]));
ibuf N51P_1_2 (.o(FF_LA[1]), .i(XFF_LA[1]));
ibuf N51P_1_1 (.o(FF_LA[0]), .i(XFF_LA[0]));
obuf N50P_1_7 (.i(ERR[6]), .o(XERR[6]));
obuf N50P_1_6 (.o(XERR[5]), .i(ERR[5]));
obuf N50P_1_5 (.o(XERR[4]), .i(ERR[4]));
obuf N50P_1_4 (.o(XERR[3]), .i(ERR[3]));
obuf N50P_1_3 (.o(XERR[2]), .i(ERR[2]));
obuf N50P_1_2 (.o(XERR[1]), .i(ERR[1]));
obuf N50P_1_1 (.o(XERR[0]), .i(ERR[0]));
obuf N71P_1_5 (.i(UN_1_IBUF_67P_O[4]), .o(SPARES[4]));
obuf N71P_1_4 (.o(SPARES[3]), .i(UN_1_IBUF_67P_O[3]));
obuf N71P_1_3 (.o(SPARES[2]), .i(UN_1_IBUF_67P_O[2]));
obuf N71P_1_2 (.o(SPARES[1]), .i(UN_1_IBUF_67P_O[1]));
obuf N71P_1_1 (.o(SPARES[0]), .i(UN_1_IBUF_67P_O[0]));
obuf N75P_1 (.i(XVDD), .o(M2));
obuf N72P_1 (.i(UN_1_IBUF_68P_O), .o(SDOUT));
obuf N64P_1 (.i(UN_1_OBUF_64P_I), .o(DUMMY_OUT));
obuf N61P_1 (.i(SPECIAL_RAW), .o(xspecial_raw));
obuf N9P_1 (.i(SYNCLR24), .o(XSYNCLR24));
obuf N45P_1 (.i(gclk), .o(XGCLK));
obuf N44P_1 (.i(CLK_SYNC10), .o(XCLK_SYNC10));
obuf N43P_1 (.i(LOAD_SYNC10_n), .o(XLOAD_SYNC10_n));
obuf N42P_1 (.i(LOAD_SYNC50_n), .o(XLOAD_SYNC50_n));
obuf N41P_1 (.i(GTCLK16), .o(XGTCLK16));
obuf N40P_1 (.i(GTLOAD16_n), .o(XGTLOAD16_n));
obuf N39P_1 (.i(GTCLK24), .o(XGTCLK24));
obuf N11P_1 (.i(GTLOAD24_n), .o(XGTLOAD24_n));
obuf N10P_1 (.i(SYNCLR), .o(xsynclr));
endmodule
`uselib

module xcountsync_globals();

wire GR;
endmodule

