/* program xnf2cds.exe version EXP Tue Nov 1 11:40:30 PST 1994 (cds9174) */
/* Created from gt_countert.xcd on Wed Oct 23 11:03:11 1996 */
/* PART 3030PC44-100 */

`timescale 1 ns/100 ps
`uselib dir=/cad/9404_4/share/library/xilinx/verilog3000 libext=.v
module gt_countert
(OSPARE2, OSPARE1, M2, ISPARE2, ISPARE1, RESET_n, ES24_MEMD, ES_MEMD, DOUT, DIN, BWRFLG_MEMD15, BSYNCLR24_n, BSYNCLR_n, BGTRIG_n, BFECBUSY, BERR_SYNCLR24, BERR_SYNCLR, BERR_RESET, BENW3_n, BENW1_n, BCLK, BCGTHACK2, BCGTHACK1, BCCLR_n, BBD_CGT_HI, PWRDWN_n, RDATA_n, RTRIG, P20, PROGRAM_n, CCLK, P43, P44);
   output OSPARE2;
   output OSPARE1;
   output M2;
   input ISPARE2;
   input ISPARE1;
   input RESET_n;
   inout ES24_MEMD;
   inout ES_MEMD;
   output DOUT;
   input DIN;
   input BWRFLG_MEMD15;
   input BSYNCLR24_n;
   input BSYNCLR_n;
   input BGTRIG_n;
   input BFECBUSY;
   output BERR_SYNCLR24;
   output BERR_SYNCLR;
   input BERR_RESET;
   input BENW3_n;
   input BENW1_n;
   input BCLK;
   input BCGTHACK2;
   input BCGTHACK1;
   input BCCLR_n;
   inout [7:0] BBD_CGT_HI;
   input PWRDWN_n;
   output RDATA_n;
   input RTRIG;
   inout P20;
   input PROGRAM_n;
   input CCLK;
   inout P43;
   inout P44;
wire [0:0] N26P_2_I47;
wire [0:0] N25P_2_I47;
wire [0:0] N24P_2_I47;
wire [7:0] N18P_4_M1;
wire [7:0] N18P_4_M0;
wire [0:0] N7P_1_I57_1_TQ;
wire [0:0] N7P_1_I52_1_TQ;
wire [0:0] N7P_1_I51_1_TQ;
wire [0:0] N7P_1_I48_1_TQ;
wire [0:0] N7P_1_I45_1_TQ;
wire [0:0] N7P_1_I43_1_TQ;
wire [0:0] N7P_1_I40_1_TQ;
wire [0:0] N7P_1_I38_1_TQ;
wire [0:0] N7P_1_I37_1_TQ;
wire [0:0] N7P_1_I35_1_TQ;
wire [0:0] N7P_1_I32_1_TQ;
wire [0:0] N7P_1_I31_1_TQ;
wire [0:0] N7P_1_I30_1_TQ;
wire [0:0] N7P_1_I27_1_TQ;
wire [0:0] N7P_1_I25_1_TQ;
wire [0:0] N7P_1_I24_1_TQ;
wire [0:0] N4P_1_I34_1_TQ;
wire [0:0] N4P_1_I30_1_TQ;
wire [0:0] N4P_1_I28_1_TQ;
wire [0:0] N4P_1_I26_1_TQ;
wire [0:0] N4P_1_I23_1_TQ;
wire [0:0] N4P_1_I20_1_TQ;
wire [0:0] N4P_1_I18_1_TQ;
wire [0:0] N4P_1_I15_1_TQ;
wire [0:0] N3P_1_I44_1_TQ;
wire [0:0] N3P_1_I44_1_MD;
wire [0:0] N3P_1_I44_1_I8_1_M1;
wire [0:0] N3P_1_I44_1_I8_1_M0;
wire [0:0] N3P_1_I43_1_TQ;
wire [0:0] N3P_1_I43_1_MD;
wire [0:0] N3P_1_I43_1_I8_1_M1;
wire [0:0] N3P_1_I43_1_I8_1_M0;
wire [0:0] N3P_1_I39_1_TQ;
wire [0:0] N3P_1_I39_1_MD;
wire [0:0] N3P_1_I39_1_I8_1_M1;
wire [0:0] N3P_1_I39_1_I8_1_M0;
wire [0:0] N3P_1_I36_1_TQ;
wire [0:0] N3P_1_I36_1_MD;
wire [0:0] N3P_1_I36_1_I8_1_M1;
wire [0:0] N3P_1_I36_1_I8_1_M0;
wire [0:0] N3P_1_I35_1_TQ;
wire [0:0] N3P_1_I35_1_MD;
wire [0:0] N3P_1_I35_1_I8_1_M1;
wire [0:0] N3P_1_I35_1_I8_1_M0;
wire [0:0] N3P_1_I31_1_TQ;
wire [0:0] N3P_1_I31_1_MD;
wire [0:0] N3P_1_I31_1_I8_1_M1;
wire [0:0] N3P_1_I31_1_I8_1_M0;
wire [0:0] N3P_1_I26_1_TQ;
wire [0:0] N3P_1_I26_1_MD;
wire [0:0] N3P_1_I26_1_I8_1_M1;
wire [0:0] N3P_1_I26_1_I8_1_M0;
wire [0:0] N3P_1_I25_1_TQ;
wire [0:0] N3P_1_I25_1_MD;
wire [0:0] N3P_1_I25_1_I8_1_M1;
wire [0:0] N3P_1_I25_1_I8_1_M0;
wire [7:0] UN_1_BUFE8_39P_O;
wire [7:0] CGT_HIM1;
wire [7:0] CGT_HI;
wire [15:0] CGT;
wire [7:0] BD2_CGT_HI;
wire [7:0] BD1_CGT_HI;
wire [7:0] BD_CGT_HI;
supply1 XVDD;
supply0 XGND;

parameter SDFFILE = "/tape/snopcb/vdwater/fec32/gtcounter/gt_countert/verilog_lib/gt_countert.sdf";
parameter SDFCONFIG = "___unspecified___";

initial $sdf_annotate(SDFFILE);

and2b1 N18P_4_I7_1_8 (.i0(UN_4_AND2_35P_O), .o(N18P_4_M0[7]), .i1(BD1_CGT_HI[7]));
and2b1 N18P_4_I7_1_7 (.i1(BD1_CGT_HI[6]), .o(N18P_4_M0[6]), .i0(UN_4_AND2_35P_O));
and2b1 N18P_4_I7_1_6 (.i1(BD1_CGT_HI[5]), .o(N18P_4_M0[5]), .i0(UN_4_AND2_35P_O));
and2b1 N18P_4_I7_1_5 (.i1(BD1_CGT_HI[4]), .o(N18P_4_M0[4]), .i0(UN_4_AND2_35P_O));
and2b1 N18P_4_I7_1_4 (.i1(BD1_CGT_HI[3]), .o(N18P_4_M0[3]), .i0(UN_4_AND2_35P_O));
and2b1 N18P_4_I7_1_3 (.i1(BD1_CGT_HI[2]), .o(N18P_4_M0[2]), .i0(UN_4_AND2_35P_O));
and2b1 N18P_4_I7_1_2 (.i1(BD1_CGT_HI[1]), .o(N18P_4_M0[1]), .i0(UN_4_AND2_35P_O));
and2b1 N18P_4_I7_1_1 (.i1(BD1_CGT_HI[0]), .o(N18P_4_M0[0]), .i0(UN_4_AND2_35P_O));
or2 N18P_4_I5_1_8 (.i0(N18P_4_M1[7]), .o(BD_CGT_HI[7]), .i1(N18P_4_M0[7]));
or2 N18P_4_I5_1_7 (.i1(N18P_4_M0[6]), .o(BD_CGT_HI[6]), .i0(N18P_4_M1[6]));
or2 N18P_4_I5_1_6 (.i1(N18P_4_M0[5]), .o(BD_CGT_HI[5]), .i0(N18P_4_M1[5]));
or2 N18P_4_I5_1_5 (.i1(N18P_4_M0[4]), .o(BD_CGT_HI[4]), .i0(N18P_4_M1[4]));
or2 N18P_4_I5_1_4 (.i1(N18P_4_M0[3]), .o(BD_CGT_HI[3]), .i0(N18P_4_M1[3]));
or2 N18P_4_I5_1_3 (.i1(N18P_4_M0[2]), .o(BD_CGT_HI[2]), .i0(N18P_4_M1[2]));
or2 N18P_4_I5_1_2 (.i1(N18P_4_M0[1]), .o(BD_CGT_HI[1]), .i0(N18P_4_M1[1]));
or2 N18P_4_I5_1_1 (.i1(N18P_4_M0[0]), .o(BD_CGT_HI[0]), .i0(N18P_4_M1[0]));
and2 N18P_4_I6_1_8 (.i0(BD2_CGT_HI[7]), .o(N18P_4_M1[7]), .i1(UN_4_AND2_35P_O));
and2 N18P_4_I6_1_7 (.i1(UN_4_AND2_35P_O), .o(N18P_4_M1[6]), .i0(BD2_CGT_HI[6]));
and2 N18P_4_I6_1_6 (.i1(UN_4_AND2_35P_O), .o(N18P_4_M1[5]), .i0(BD2_CGT_HI[5]));
and2 N18P_4_I6_1_5 (.i1(UN_4_AND2_35P_O), .o(N18P_4_M1[4]), .i0(BD2_CGT_HI[4]));
and2 N18P_4_I6_1_4 (.i1(UN_4_AND2_35P_O), .o(N18P_4_M1[3]), .i0(BD2_CGT_HI[3]));
and2 N18P_4_I6_1_3 (.i1(UN_4_AND2_35P_O), .o(N18P_4_M1[2]), .i0(BD2_CGT_HI[2]));
and2 N18P_4_I6_1_2 (.i1(UN_4_AND2_35P_O), .o(N18P_4_M1[1]), .i0(BD2_CGT_HI[1]));
and2 N18P_4_I6_1_1 (.i1(UN_4_AND2_35P_O), .o(N18P_4_M1[0]), .i0(BD2_CGT_HI[0]));
fdce N11P_4_I19_1 (.q(UN_4_OBUFE_87P_I), .d(BD_CGT_HI[3]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
fdce N11P_4_I22_1 (.q(UN_4_OBUFE_84P_I), .d(BD_CGT_HI[0]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
fdce N11P_4_I21_1 (.q(UN_4_OBUFE_88P_I), .d(BD_CGT_HI[4]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
fdce N11P_4_I20_1 (.q(UN_4_OBUFE_89P_I), .d(BD_CGT_HI[5]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
fdce N11P_4_I27_1 (.q(UN_4_OBUFE_85P_I), .d(BD_CGT_HI[1]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
fdce N11P_4_I26_1 (.q(UN_4_OBUFE_90P_I), .d(BD_CGT_HI[6]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
fdce N11P_4_I29_1 (.q(UN_4_OBUFE_91P_I), .d(BD_CGT_HI[7]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
fdce N11P_4_I24_1 (.q(UN_4_OBUFE_86P_I), .d(BD_CGT_HI[2]), .ce(N11P_4_GB), .c(ENWRITE1_n), .clr(XGND), .gr(RESET_n));
inv N11P_4_I23_1 (.i(UN_4_NOR2_36P_O), .o(N11P_4_GB));
obuft N90P_4_I5_1 (.i(UN_4_OBUFE_90P_I), .o(BBD_CGT_HI[6]), .t(N90P_4_T));
inv N90P_4_I4_1 (.i(ENWRITE3), .o(N90P_4_T));
obuft N89P_4_I5_1 (.i(UN_4_OBUFE_89P_I), .o(BBD_CGT_HI[5]), .t(N89P_4_T));
inv N89P_4_I4_1 (.i(ENWRITE3), .o(N89P_4_T));
obuft N88P_4_I5_1 (.i(UN_4_OBUFE_88P_I), .o(BBD_CGT_HI[4]), .t(N88P_4_T));
inv N88P_4_I4_1 (.i(ENWRITE3), .o(N88P_4_T));
obuft N87P_4_I5_1 (.i(UN_4_OBUFE_87P_I), .o(BBD_CGT_HI[3]), .t(N87P_4_T));
inv N87P_4_I4_1 (.i(ENWRITE3), .o(N87P_4_T));
obuft N86P_4_I5_1 (.i(UN_4_OBUFE_86P_I), .o(BBD_CGT_HI[2]), .t(N86P_4_T));
inv N86P_4_I4_1 (.i(ENWRITE3), .o(N86P_4_T));
obuft N84P_4_I5_1 (.i(UN_4_OBUFE_84P_I), .o(BBD_CGT_HI[0]), .t(N84P_4_T));
inv N84P_4_I4_1 (.i(ENWRITE3), .o(N84P_4_T));
obuft N70P_4_I5_1 (.i(UN_4_FDC_69P_Q), .o(ES24_MEMD), .t(N70P_4_T));
inv N70P_4_I4_1 (.i(ENWRITE1), .o(N70P_4_T));
obuft N66P_4_I5_1 (.i(UN_4_FDC_20P_Q), .o(ES_MEMD), .t(N66P_4_T));
inv N66P_4_I4_1 (.i(ENWRITE1), .o(N66P_4_T));
obuft N91P_4_I5_1 (.i(UN_4_OBUFE_91P_I), .o(BBD_CGT_HI[7]), .t(N91P_4_T));
inv N91P_4_I4_1 (.i(ENWRITE3), .o(N91P_4_T));
obuft N85P_4_I5_1 (.i(UN_4_OBUFE_85P_I), .o(BBD_CGT_HI[1]), .t(N85P_4_T));
inv N85P_4_I4_1 (.i(ENWRITE3), .o(N85P_4_T));
and4 N81P_3_I56_1 (.i3(N81P_3_AB03), .i2(N81P_3_AB47), .i0(N81P_3_ABCF), .o(ENCCLR), .i1(N81P_3_AB8B));
and4 N81P_3_I53_1 (.i3(N81P_3_AB4), .i2(N81P_3_AB5), .i0(N81P_3_AB7), .o(N81P_3_AB47), .i1(N81P_3_AB6));
and4 N81P_3_I49_1 (.i3(N81P_3_AB0), .i2(N81P_3_AB1), .i0(N81P_3_AB3), .o(N81P_3_AB03), .i1(N81P_3_AB2));
and4 N81P_3_I41_1 (.i3(N81P_3_AB12), .i2(N81P_3_AB13), .i0(N81P_3_AB15), .o(N81P_3_ABCF), .i1(N81P_3_AB14));
and4 N81P_3_I40_1 (.i3(N81P_3_AB8), .i2(N81P_3_AB9), .i0(N81P_3_AB11), .o(N81P_3_AB8B), .i1(N81P_3_AB10));
xnor2 N81P_3_I55_1 (.i0(XVDD), .o(N81P_3_AB1), .i1(CGT[1]));
xnor2 N81P_3_I54_1 (.i0(XVDD), .o(N81P_3_AB13), .i1(CGT[13]));
xnor2 N81P_3_I46_1 (.i0(XVDD), .o(N81P_3_AB2), .i1(CGT[2]));
xnor2 N81P_3_I42_1 (.i0(XVDD), .o(N81P_3_AB6), .i1(CGT[6]));
xnor2 N81P_3_I47_1 (.i0(XVDD), .o(N81P_3_AB4), .i1(CGT[4]));
xnor2 N81P_3_I58_1 (.i0(XVDD), .o(N81P_3_AB10), .i1(CGT[10]));
xnor2 N81P_3_I57_1 (.i0(XGND), .o(N81P_3_AB15), .i1(CGT[15]));
xnor2 N81P_3_I52_1 (.i0(XVDD), .o(N81P_3_AB12), .i1(CGT[12]));
xnor2 N81P_3_I51_1 (.i0(XVDD), .o(N81P_3_AB5), .i1(CGT[5]));
xnor2 N81P_3_I45_1 (.i0(XVDD), .o(N81P_3_AB7), .i1(CGT[7]));
xnor2 N81P_3_I44_1 (.i0(XVDD), .o(N81P_3_AB0), .i1(CGT[0]));
xnor2 N81P_3_I43_1 (.i0(XVDD), .o(N81P_3_AB11), .i1(CGT[11]));
xnor2 N81P_3_I39_1 (.i0(XVDD), .o(N81P_3_AB9), .i1(CGT[9]));
xnor2 N81P_3_I38_1 (.i0(XVDD), .o(N81P_3_AB3), .i1(CGT[3]));
xnor2 N81P_3_I37_1 (.i0(XVDD), .o(N81P_3_AB14), .i1(CGT[14]));
xnor2 N81P_3_I36_1 (.i0(XVDD), .o(N81P_3_AB8), .i1(CGT[8]));
nand5 N26P_2_I10_1 (.i4(N26P_2_I47[0]), .i3(CGT_HI[3]), .i2(CGT_HI[2]), .i0(CGT_HI[0]), .o(UN_2_AND2_1P_I0), .i1(CGT_HI[1]));
and4 N26P_2_I12_1 (.i3(CGT_HI[7]), .i2(CGT_HI[6]), .i0(CGT_HI[4]), .o(N26P_2_I47[0]), .i1(CGT_HI[5]));
nand5 N25P_2_I10_1 (.i4(N25P_2_I47[0]), .i3(CGT[11]), .i2(CGT[10]), .i0(CGT[8]), .o(UN_2_NAND8_25P_O), .i1(CGT[9]));
and4 N25P_2_I12_1 (.i3(CGT[15]), .i2(CGT[14]), .i0(CGT[12]), .o(N25P_2_I47[0]), .i1(CGT[13]));
nand5 N24P_2_I10_1 (.i4(N24P_2_I47[0]), .i3(CGT[3]), .i2(CGT[2]), .i0(CGT[0]), .o(UN_2_NAND8_24P_O), .i1(CGT[1]));
and4 N24P_2_I12_1 (.i3(CGT[7]), .i2(CGT[6]), .i0(CGT[4]), .o(N24P_2_I47[0]), .i1(CGT[5]));
fdce N7P_1_I57_1_I7_1 (.q(CGT[5]), .d(N7P_1_I57_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I57_1_I8_1 (.i0(N7P_1_T5), .o(N7P_1_I57_1_TQ[0]), .i1(CGT[5]));
fdce N7P_1_I52_1_I7_1 (.q(CGT[0]), .d(N7P_1_I52_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I52_1_I8_1 (.i0(XVDD), .o(N7P_1_I52_1_TQ[0]), .i1(CGT[0]));
fdce N7P_1_I51_1_I7_1 (.q(CGT[12]), .d(N7P_1_I51_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I51_1_I8_1 (.i0(N7P_1_T12), .o(N7P_1_I51_1_TQ[0]), .i1(CGT[12]));
fdce N7P_1_I48_1_I7_1 (.q(CGT[13]), .d(N7P_1_I48_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I48_1_I8_1 (.i0(N7P_1_T13), .o(N7P_1_I48_1_TQ[0]), .i1(CGT[13]));
fdce N7P_1_I45_1_I7_1 (.q(CGT[10]), .d(N7P_1_I45_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I45_1_I8_1 (.i0(N7P_1_T10), .o(N7P_1_I45_1_TQ[0]), .i1(CGT[10]));
fdce N7P_1_I40_1_I7_1 (.q(CGT[14]), .d(N7P_1_I40_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I40_1_I8_1 (.i0(N7P_1_T14), .o(N7P_1_I40_1_TQ[0]), .i1(CGT[14]));
fdce N7P_1_I43_1_I7_1 (.q(CGT[8]), .d(N7P_1_I43_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I43_1_I8_1 (.i0(N7P_1_T8), .o(N7P_1_I43_1_TQ[0]), .i1(CGT[8]));
fdce N7P_1_I38_1_I7_1 (.q(CGT[4]), .d(N7P_1_I38_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I38_1_I8_1 (.i0(N7P_1_T4), .o(N7P_1_I38_1_TQ[0]), .i1(CGT[4]));
fdce N7P_1_I32_1_I7_1 (.q(CGT[2]), .d(N7P_1_I32_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I32_1_I8_1 (.i0(N7P_1_T2), .o(N7P_1_I32_1_TQ[0]), .i1(CGT[2]));
fdce N7P_1_I27_1_I7_1 (.q(CGT[1]), .d(N7P_1_I27_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I27_1_I8_1 (.i0(CGT[0]), .o(N7P_1_I27_1_TQ[0]), .i1(CGT[1]));
fdce N7P_1_I25_1_I7_1 (.q(CGT[7]), .d(N7P_1_I25_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I25_1_I8_1 (.i0(N7P_1_T7), .o(N7P_1_I25_1_TQ[0]), .i1(CGT[7]));
fdce N7P_1_I37_1_I7_1 (.q(CGT[9]), .d(N7P_1_I37_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I37_1_I8_1 (.i0(N7P_1_T9), .o(N7P_1_I37_1_TQ[0]), .i1(CGT[9]));
fdce N7P_1_I35_1_I7_1 (.q(CGT[6]), .d(N7P_1_I35_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I35_1_I8_1 (.i0(N7P_1_T6), .o(N7P_1_I35_1_TQ[0]), .i1(CGT[6]));
fdce N7P_1_I31_1_I7_1 (.q(CGT[11]), .d(N7P_1_I31_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I31_1_I8_1 (.i0(N7P_1_T11), .o(N7P_1_I31_1_TQ[0]), .i1(CGT[11]));
fdce N7P_1_I30_1_I7_1 (.q(CGT[3]), .d(N7P_1_I30_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I30_1_I8_1 (.i0(N7P_1_T3), .o(N7P_1_I30_1_TQ[0]), .i1(CGT[3]));
fdce N7P_1_I24_1_I7_1 (.q(CGT[15]), .d(N7P_1_I24_1_TQ[0]), .ce(XVDD), .c(LOWINC), .clr(UN_1_CB16CE_7P_CLR), .gr(RESET_n));
xor2 N7P_1_I24_1_I8_1 (.i0(N7P_1_T15), .o(N7P_1_I24_1_TQ[0]), .i1(CGT[15]));
and3 N7P_1_I72_1 (.i2(CGT[0]), .i0(CGT[2]), .o(N7P_1_T3), .i1(CGT[1]));
and3 N7P_1_I70_1 (.i2(N7P_1_T8), .i0(CGT[9]), .o(N7P_1_T10), .i1(CGT[8]));
and3 N7P_1_I64_1 (.i2(N7P_1_T12), .i0(CGT[13]), .o(N7P_1_T14), .i1(CGT[12]));
and3 N7P_1_I61_1 (.i2(N7P_1_T4), .i0(CGT[5]), .o(N7P_1_T6), .i1(CGT[4]));
and5 N7P_1_I73_1 (.i4(N7P_1_T12), .i3(CGT[12]), .i2(CGT[13]), .i0(CGT[15]), .o(N7P_1_TC), .i1(CGT[14]));
and5 N7P_1_I66_1 (.i4(N7P_1_T8), .i3(CGT[8]), .i2(CGT[9]), .i0(CGT[11]), .o(N7P_1_T12), .i1(CGT[10]));
and5 N7P_1_I63_1 (.i4(N7P_1_T4), .i3(CGT[4]), .i2(CGT[5]), .i0(CGT[7]), .o(N7P_1_T8), .i1(CGT[6]));
and4 N7P_1_I74_1 (.i3(N7P_1_T12), .i2(CGT[12]), .i0(CGT[14]), .o(N7P_1_T15), .i1(CGT[13]));
and4 N7P_1_I67_1 (.i3(N7P_1_T4), .i2(CGT[4]), .i0(CGT[6]), .o(N7P_1_T7), .i1(CGT[5]));
and4 N7P_1_I62_1 (.i3(CGT[0]), .i2(CGT[1]), .i0(CGT[3]), .o(N7P_1_T4), .i1(CGT[2]));
and4 N7P_1_I59_1 (.i3(N7P_1_T8), .i2(CGT[8]), .i0(CGT[10]), .o(N7P_1_T11), .i1(CGT[9]));
and2 N7P_1_I69_1 (.i0(CGT[4]), .o(N7P_1_T5), .i1(N7P_1_T4));
and2 N7P_1_I68_1 (.i0(CGT[8]), .o(N7P_1_T9), .i1(N7P_1_T8));
and2 N7P_1_I65_1 (.i0(XVDD), .o(N7P_1_CEO), .i1(N7P_1_TC));
and2 N7P_1_I60_1 (.i0(CGT[1]), .o(N7P_1_T2), .i1(CGT[0]));
and2 N7P_1_I58_1 (.i0(CGT[12]), .o(N7P_1_T13), .i1(N7P_1_T12));
fdce N4P_1_I23_1_I7_1 (.q(CGT_HI[5]), .d(N4P_1_I23_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I23_1_I8_1 (.i0(N4P_1_T5), .o(N4P_1_I23_1_TQ[0]), .i1(CGT_HI[5]));
fdce N4P_1_I20_1_I7_1 (.q(CGT_HI[2]), .d(N4P_1_I20_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I20_1_I8_1 (.i0(N4P_1_T2), .o(N4P_1_I20_1_TQ[0]), .i1(CGT_HI[2]));
fdce N4P_1_I18_1_I7_1 (.q(CGT_HI[3]), .d(N4P_1_I18_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I18_1_I8_1 (.i0(N4P_1_T3), .o(N4P_1_I18_1_TQ[0]), .i1(CGT_HI[3]));
fdce N4P_1_I15_1_I7_1 (.q(CGT_HI[7]), .d(N4P_1_I15_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I15_1_I8_1 (.i0(N4P_1_T7), .o(N4P_1_I15_1_TQ[0]), .i1(CGT_HI[7]));
fdce N4P_1_I26_1_I7_1 (.q(CGT_HI[1]), .d(N4P_1_I26_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I26_1_I8_1 (.i0(CGT_HI[0]), .o(N4P_1_I26_1_TQ[0]), .i1(CGT_HI[1]));
fdce N4P_1_I34_1_I7_1 (.q(CGT_HI[0]), .d(N4P_1_I34_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I34_1_I8_1 (.i0(XVDD), .o(N4P_1_I34_1_TQ[0]), .i1(CGT_HI[0]));
fdce N4P_1_I30_1_I7_1 (.q(CGT_HI[4]), .d(N4P_1_I30_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I30_1_I8_1 (.i0(N4P_1_T4), .o(N4P_1_I30_1_TQ[0]), .i1(CGT_HI[4]));
fdce N4P_1_I28_1_I7_1 (.q(CGT_HI[6]), .d(N4P_1_I28_1_TQ[0]), .ce(XVDD), .c(UPINC), .clr(UN_1_CB8CE_4P_CLR), .gr(RESET_n));
xor2 N4P_1_I28_1_I8_1 (.i0(N4P_1_T6), .o(N4P_1_I28_1_TQ[0]), .i1(CGT_HI[6]));
and3 N4P_1_I32_1 (.i2(CGT_HI[0]), .i0(CGT_HI[2]), .o(N4P_1_T3), .i1(CGT_HI[1]));
and3 N4P_1_I33_1 (.i2(N4P_1_T4), .i0(CGT_HI[5]), .o(N4P_1_T6), .i1(CGT_HI[4]));
and5 N4P_1_I25_1 (.i4(N4P_1_T4), .i3(CGT_HI[4]), .i2(CGT_HI[5]), .i0(CGT_HI[7]), .o(N4P_1_TC), .i1(CGT_HI[6]));
and4 N4P_1_I16_1 (.i3(CGT_HI[0]), .i2(CGT_HI[1]), .i0(CGT_HI[3]), .o(N4P_1_T4), .i1(CGT_HI[2]));
and4 N4P_1_I24_1 (.i3(N4P_1_T4), .i2(CGT_HI[4]), .i0(CGT_HI[6]), .o(N4P_1_T7), .i1(CGT_HI[5]));
and2 N4P_1_I22_1 (.i0(XVDD), .o(N4P_1_CEO), .i1(N4P_1_TC));
and2 N4P_1_I21_1 (.i0(CGT_HI[4]), .o(N4P_1_T5), .i1(N4P_1_T4));
and2 N4P_1_I29_1 (.i0(CGT_HI[1]), .o(N4P_1_T2), .i1(CGT_HI[0]));
and2b1 N3P_1_I44_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I44_1_I8_1_M0[0]), .i1(N3P_1_I44_1_TQ[0]));
or2 N3P_1_I44_1_I8_1_I5_1 (.i0(N3P_1_I44_1_I8_1_M1[0]), .o(N3P_1_I44_1_MD[0]), .i1(N3P_1_I44_1_I8_1_M0[0]));
and2 N3P_1_I44_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[6]), .o(N3P_1_I44_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I44_1_I12_1 (.q(CGT_HIM1[6]), .d(N3P_1_I44_1_MD[0]), .ce(N3P_1_I44_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I44_1_I13_1 (.i0(XVDD), .o(N3P_1_I44_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I44_1_I9_1 (.i0(N3P_1_T6), .o(N3P_1_I44_1_TQ[0]), .i1(CGT_HIM1[6]));
and2b1 N3P_1_I43_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I43_1_I8_1_M0[0]), .i1(N3P_1_I43_1_TQ[0]));
or2 N3P_1_I43_1_I8_1_I5_1 (.i0(N3P_1_I43_1_I8_1_M1[0]), .o(N3P_1_I43_1_MD[0]), .i1(N3P_1_I43_1_I8_1_M0[0]));
and2 N3P_1_I43_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[5]), .o(N3P_1_I43_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I43_1_I12_1 (.q(CGT_HIM1[5]), .d(N3P_1_I43_1_MD[0]), .ce(N3P_1_I43_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I43_1_I13_1 (.i0(XVDD), .o(N3P_1_I43_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I43_1_I9_1 (.i0(N3P_1_T5), .o(N3P_1_I43_1_TQ[0]), .i1(CGT_HIM1[5]));
and2b1 N3P_1_I39_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I39_1_I8_1_M0[0]), .i1(N3P_1_I39_1_TQ[0]));
or2 N3P_1_I39_1_I8_1_I5_1 (.i0(N3P_1_I39_1_I8_1_M1[0]), .o(N3P_1_I39_1_MD[0]), .i1(N3P_1_I39_1_I8_1_M0[0]));
and2 N3P_1_I39_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[7]), .o(N3P_1_I39_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I39_1_I12_1 (.q(CGT_HIM1[7]), .d(N3P_1_I39_1_MD[0]), .ce(N3P_1_I39_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I39_1_I13_1 (.i0(XVDD), .o(N3P_1_I39_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I39_1_I9_1 (.i0(N3P_1_T7), .o(N3P_1_I39_1_TQ[0]), .i1(CGT_HIM1[7]));
and2b1 N3P_1_I26_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I26_1_I8_1_M0[0]), .i1(N3P_1_I26_1_TQ[0]));
or2 N3P_1_I26_1_I8_1_I5_1 (.i0(N3P_1_I26_1_I8_1_M1[0]), .o(N3P_1_I26_1_MD[0]), .i1(N3P_1_I26_1_I8_1_M0[0]));
and2 N3P_1_I26_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[2]), .o(N3P_1_I26_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I26_1_I12_1 (.q(CGT_HIM1[2]), .d(N3P_1_I26_1_MD[0]), .ce(N3P_1_I26_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I26_1_I13_1 (.i0(XVDD), .o(N3P_1_I26_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I26_1_I9_1 (.i0(N3P_1_T2), .o(N3P_1_I26_1_TQ[0]), .i1(CGT_HIM1[2]));
and2b1 N3P_1_I25_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I25_1_I8_1_M0[0]), .i1(N3P_1_I25_1_TQ[0]));
or2 N3P_1_I25_1_I8_1_I5_1 (.i0(N3P_1_I25_1_I8_1_M1[0]), .o(N3P_1_I25_1_MD[0]), .i1(N3P_1_I25_1_I8_1_M0[0]));
and2 N3P_1_I25_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[4]), .o(N3P_1_I25_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I25_1_I12_1 (.q(CGT_HIM1[4]), .d(N3P_1_I25_1_MD[0]), .ce(N3P_1_I25_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I25_1_I13_1 (.i0(XVDD), .o(N3P_1_I25_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I25_1_I9_1 (.i0(N3P_1_T4), .o(N3P_1_I25_1_TQ[0]), .i1(CGT_HIM1[4]));
and2b1 N3P_1_I36_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I36_1_I8_1_M0[0]), .i1(N3P_1_I36_1_TQ[0]));
or2 N3P_1_I36_1_I8_1_I5_1 (.i0(N3P_1_I36_1_I8_1_M1[0]), .o(N3P_1_I36_1_MD[0]), .i1(N3P_1_I36_1_I8_1_M0[0]));
and2 N3P_1_I36_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[3]), .o(N3P_1_I36_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I36_1_I12_1 (.q(CGT_HIM1[3]), .d(N3P_1_I36_1_MD[0]), .ce(N3P_1_I36_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I36_1_I13_1 (.i0(XVDD), .o(N3P_1_I36_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I36_1_I9_1 (.i0(N3P_1_T3), .o(N3P_1_I36_1_TQ[0]), .i1(CGT_HIM1[3]));
and2b1 N3P_1_I35_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I35_1_I8_1_M0[0]), .i1(N3P_1_I35_1_TQ[0]));
or2 N3P_1_I35_1_I8_1_I5_1 (.i0(N3P_1_I35_1_I8_1_M1[0]), .o(N3P_1_I35_1_MD[0]), .i1(N3P_1_I35_1_I8_1_M0[0]));
and2 N3P_1_I35_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[0]), .o(N3P_1_I35_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I35_1_I12_1 (.q(CGT_HIM1[0]), .d(N3P_1_I35_1_MD[0]), .ce(N3P_1_I35_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I35_1_I13_1 (.i0(XVDD), .o(N3P_1_I35_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I35_1_I9_1 (.i0(XVDD), .o(N3P_1_I35_1_TQ[0]), .i1(CGT_HIM1[0]));
and2b1 N3P_1_I31_1_I8_1_I7_1 (.i0(UN_1_CB8CLE_3P_L), .o(N3P_1_I31_1_I8_1_M0[0]), .i1(N3P_1_I31_1_TQ[0]));
or2 N3P_1_I31_1_I8_1_I5_1 (.i0(N3P_1_I31_1_I8_1_M1[0]), .o(N3P_1_I31_1_MD[0]), .i1(N3P_1_I31_1_I8_1_M0[0]));
and2 N3P_1_I31_1_I8_1_I6_1 (.i0(UN_1_BUFE8_39P_O[1]), .o(N3P_1_I31_1_I8_1_M1[0]), .i1(UN_1_CB8CLE_3P_L));
fdce N3P_1_I31_1_I12_1 (.q(CGT_HIM1[1]), .d(N3P_1_I31_1_MD[0]), .ce(N3P_1_I31_1_L_CE), .c(UN_1_CB8CLE_3P_C), .clr(UN_1_AND2_95P_O), .gr(RESET_n));
or2 N3P_1_I31_1_I13_1 (.i0(XVDD), .o(N3P_1_I31_1_L_CE), .i1(UN_1_CB8CLE_3P_L));
xor2 N3P_1_I31_1_I9_1 (.i0(CGT_HIM1[0]), .o(N3P_1_I31_1_TQ[0]), .i1(CGT_HIM1[1]));
and3 N3P_1_I27_1 (.i2(N3P_1_T4), .i0(CGT_HIM1[5]), .o(N3P_1_T6), .i1(CGT_HIM1[4]));
and3 N3P_1_I29_1 (.i2(CGT_HIM1[0]), .i0(CGT_HIM1[2]), .o(N3P_1_T3), .i1(CGT_HIM1[1]));
and5 N3P_1_I37_1 (.i4(N3P_1_T4), .i3(CGT_HIM1[4]), .i2(CGT_HIM1[5]), .i0(CGT_HIM1[7]), .o(N3P_1_TC), .i1(CGT_HIM1[6]));
and4 N3P_1_I38_1 (.i3(CGT_HIM1[0]), .i2(CGT_HIM1[1]), .i0(CGT_HIM1[3]), .o(N3P_1_T4), .i1(CGT_HIM1[2]));
and4 N3P_1_I33_1 (.i3(N3P_1_T4), .i2(CGT_HIM1[4]), .i0(CGT_HIM1[6]), .o(N3P_1_T7), .i1(CGT_HIM1[5]));
and2 N3P_1_I32_1 (.i0(XVDD), .o(N3P_1_CEO), .i1(N3P_1_TC));
and2 N3P_1_I34_1 (.i0(CGT_HIM1[4]), .o(N3P_1_T5), .i1(N3P_1_T4));
and2 N3P_1_I30_1 (.i0(CGT_HIM1[1]), .o(N3P_1_T2), .i1(CGT_HIM1[0]));
buft N39P_1_I37_1 (.i(CGT_HI[0]), .o(UN_1_BUFE8_39P_O[0]), .t(N39P_1_T));
buft N39P_1_I36_1 (.i(CGT_HI[5]), .o(UN_1_BUFE8_39P_O[5]), .t(N39P_1_T));
buft N39P_1_I35_1 (.i(CGT_HI[6]), .o(UN_1_BUFE8_39P_O[6]), .t(N39P_1_T));
buft N39P_1_I34_1 (.i(CGT_HI[3]), .o(UN_1_BUFE8_39P_O[3]), .t(N39P_1_T));
buft N39P_1_I33_1 (.i(CGT_HI[7]), .o(UN_1_BUFE8_39P_O[7]), .t(N39P_1_T));
buft N39P_1_I31_1 (.i(CGT_HI[2]), .o(UN_1_BUFE8_39P_O[2]), .t(N39P_1_T));
buft N39P_1_I30_1 (.i(CGT_HI[1]), .o(UN_1_BUFE8_39P_O[1]), .t(N39P_1_T));
buft N39P_1_I28_1 (.i(CGT_HI[4]), .o(UN_1_BUFE8_39P_O[4]), .t(N39P_1_T));
inv N39P_1_I29_1 (.i(SYNCLR24_GATE), .o(N39P_1_T));
fdce N69P_4_I8_1 (.q(UN_4_FDC_69P_Q), .d(XVDD), .ce(XVDD), .c(ERR_SYNCLR24), .clr(UN_4_FDC_69P_CLR), .gr(RESET_n));
fdce N20P_4_I8_1 (.q(UN_4_FDC_20P_Q), .d(XVDD), .ce(XVDD), .c(ERR_SYNCLR), .clr(UN_4_FDC_20P_CLR), .gr(RESET_n));
fdce N38P_3_I8_1 (.q(SYNCLR24_D2), .d(SYNCLR24_D1), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
fdce N37P_3_I8_1 (.q(SYNCLR24_D1), .d(UN_3_FDC_34P_Q), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
fdce N31P_3_I8_1 (.q(UN_3_FDC_30P_D), .d(XVDD), .ce(XVDD), .c(SYNCLR_n), .clr(UN_3_FDC_31P_CLR), .gr(RESET_n));
fdce N30P_3_I8_1 (.q(SYNCLR_D1), .d(UN_3_FDC_30P_D), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
fdce N29P_3_I8_1 (.q(SYNCLR_D2), .d(SYNCLR_D1), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
fdce N111P_3_I8_1 (.q(UN_3_FDC_109P_D), .d(XVDD), .ce(XVDD), .c(ENWRITE1_n), .clr(UN_3_FDC_111P_CLR), .gr(RESET_n));
fdce N109P_3_I8_1 (.q(ENWRITE1_D1), .d(UN_3_FDC_109P_D), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
fdce N34P_3_I8_1 (.q(UN_3_FDC_34P_Q), .d(XVDD), .ce(XVDD), .c(SYNCLR24_n), .clr(UN_3_FDC_34P_CLR), .gr(RESET_n));
fdce N112P_3_I8_1 (.q(UN_3_FDC_112P_Q), .d(ENWRITE1_D1), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
fdce N47P_2_I8_1 (.q(SYNCLR24_GATE), .d(XVDD), .ce(XVDD), .c(SYNCLR24), .clr(UN_2_FDC_47P_CLR), .gr(RESET_n));
fdce N46P_2_I8_1 (.q(SYNCLR_GATE), .d(XVDD), .ce(XVDD), .c(SYNCLR), .clr(UN_2_FDC_46P_CLR), .gr(RESET_n));
fdce N40P_2_I8_1 (.q(ERR_SYNCLR24), .d(XVDD), .ce(XVDD), .c(UN_2_AND2_1P_O), .clr(UN_2_FDC_40P_CLR), .gr(RESET_n));
fdce N39P_2_I8_1 (.q(ERR_SYNCLR), .d(XVDD), .ce(XVDD), .c(UN_2_AND2_6P_O), .clr(UN_2_FDC_39P_CLR), .gr(RESET_n));
fdce N96P_1_I8_1 (.q(ENWRGT), .d(XVDD), .ce(XVDD), .c(UN_1_AND2_50P_O), .clr(UN_1_FDC_96P_CLR), .gr(RESET_n));
fdce N85P_1_I8_1 (.q(UN_1_AND2_95P_I0), .d(XVDD), .ce(XVDD), .c(SYNCLR24_D2), .clr(UN_1_FDC_85P_CLR), .gr(RESET_n));
fdce N82P_1_I8_1 (.q(UN_1_AND2_50P_I1), .d(XVDD), .ce(XVDD), .c(SYNCLR), .clr(UN_1_FDC_82P_CLR), .gr(RESET_n));
fdce N119P_1_I8_1 (.q(UN_1_FDC_118P_D), .d(XVDD), .ce(XVDD), .c(UN_1_AND2_95P_O), .clr(UN_1_FDC_119P_CLR), .gr(RESET_n));
fdce N118P_1_I8_1 (.q(UN_1_FDC_117P_D), .d(UN_1_FDC_118P_D), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
fdce N117P_1_I8_1 (.q(UN_1_FDC_117P_Q), .d(UN_1_FDC_117P_D), .ce(XVDD), .c(CLK), .clr(CCLR), .gr(RESET_n));
nor2 N36P_4 (.i0(ENREG2), .o(UN_4_NOR2_36P_O), .i1(ENREG1));
or4 N68P_4 (.i3(CCLR), .i2(ERR_RESET), .i0(ENWRITE1_D1), .o(UN_4_FDC_69P_CLR), .i1(SYNCLR24));
or4 N65P_4 (.i3(CCLR), .i2(ERR_RESET), .i0(ENWRITE1_D1), .o(UN_4_FDC_20P_CLR), .i1(SYNCLR));
obuf N2P_5 (.i(SDOUT), .o(DOUT));
obuf N3P_5 (.i(XVDD), .o(M2));
obuf N37P_4 (.i(OSP2), .o(OSPARE2));
obuf N39P_4 (.i(OSP1), .o(OSPARE1));
obuf N107P_3 (.i(ERR_SYNCLR), .o(BERR_SYNCLR));
obuf N105P_3 (.i(ERR_SYNCLR24), .o(BERR_SYNCLR24));
or3 N35P_2 (.i2(CCLR), .i0(SYNCLR), .o(UN_2_FDC_39P_CLR), .i1(ERR_RESET));
or3 N34P_2 (.i2(CCLR), .i0(SYNCLR24), .o(UN_2_FDC_40P_CLR), .i1(ERR_RESET));
ibuf N4P_5 (.i(DIN), .o(SDIN));
ibuf N57P_3 (.i(BENW1_n), .o(ENWRITE1_n));
ibuf N80P_4 (.i(BCGTHACK2), .o(CGTHACK2));
ibuf N81P_4 (.i(BCGTHACK1), .o(CGTHACK1));
ibuf N42P_4 (.i(ISPARE1), .o(ISP1));
ibuf N41P_4 (.i(ISPARE2), .o(ISP2));
ibuf N59P_3 (.i(BGTRIG_n), .o(UN_3_IBUF_59P_O));
ibuf N42P_3 (.i(BSYNCLR_n), .o(SYNCLR_n));
ibuf N114P_3 (.i(BWRFLG_MEMD15), .o(WRFLG_MEMD15));
ibuf N49P_3 (.i(BCCLR_n), .o(UN_3_IBUF_49P_O));
ibuf N46P_3 (.i(BSYNCLR24_n), .o(SYNCLR24_n));
ibuf N44P_3 (.i(BFECBUSY), .o(UN_3_IBUF_44P_O));
ibuf N43P_3 (.i(BERR_RESET), .o(ERR_RESET));
ibuf N35P_3 (.i(BCLK), .o(CLK));
ibuf N53P_3 (.i(BENW3_n), .o(UN_3_IBUF_53P_O));
pullup1 N40P_1_8 (.o(UN_1_BUFE8_39P_O[7]));
pullup1 N40P_1_7 (.o(UN_1_BUFE8_39P_O[6]));
pullup1 N40P_1_6 (.o(UN_1_BUFE8_39P_O[5]));
pullup1 N40P_1_5 (.o(UN_1_BUFE8_39P_O[4]));
pullup1 N40P_1_4 (.o(UN_1_BUFE8_39P_O[3]));
pullup1 N40P_1_3 (.o(UN_1_BUFE8_39P_O[2]));
pullup1 N40P_1_2 (.o(UN_1_BUFE8_39P_O[1]));
pullup1 N40P_1_1 (.o(UN_1_BUFE8_39P_O[0]));
or2 N110P_3 (.i0(UN_3_FDC_112P_Q), .o(UN_3_FDC_111P_CLR), .i1(CCLR));
or2 N100P_3 (.i0(SYNCLR_D2), .o(UN_3_FDC_31P_CLR), .i1(CCLR));
or2 N102P_3 (.i0(SYNCLR24_D2), .o(UN_3_FDC_34P_CLR), .i1(CCLR));
or2 N49P_2 (.i0(UN_2_NAND8_24P_O), .o(UN_2_AND2_6P_I0), .i1(UN_2_NAND8_25P_O));
or2 N48P_2 (.i0(SYNCLR24_D2), .o(UN_2_FDC_47P_CLR), .i1(CCLR));
or2 N45P_2 (.i0(SYNCLR_D2), .o(UN_2_FDC_46P_CLR), .i1(CCLR));
or2 N97P_1 (.i0(CCLR), .o(UN_1_FDC_96P_CLR), .i1(FECBUSY_n));
or2 N91P_1 (.i0(UN_1_INV_94P_O), .o(UN_1_CB8CLE_3P_C), .i1(UPINC));
or2 N77P_1 (.i0(UN_1_FDC_117P_Q), .o(UN_1_FDC_85P_CLR), .i1(CCLR));
or2 N74P_1 (.i0(UN_1_AND2_112P_O), .o(UN_1_CB8CLE_3P_L), .i1(CCLR));
or2 N73P_1 (.i0(UN_1_OR2_6P_O), .o(UN_1_CB16CE_7P_CLR), .i1(CCLR));
or2 N72P_1 (.i0(SYNCLR24_D2), .o(UN_1_CB8CE_4P_CLR), .i1(CCLR));
or2 N71P_1 (.i0(CCLR), .o(UN_1_FDC_82P_CLR), .i1(ENCCLR));
or2 N6P_1 (.i0(SYNCLR24_D2), .o(UN_1_OR2_6P_O), .i1(SYNCLR_D2));
or2 N116P_1 (.i0(UN_1_FDC_117P_Q), .o(UN_1_FDC_119P_CLR), .i1(CCLR));
xor2 N98P_1 (.i0(SYNCLR24), .o(UN_1_AND2_100P_I1), .i1(SYNCLR));
xor2 N113P_1 (.i0(SYNCLR), .o(UN_1_AND2_115P_I1), .i1(GTRIG));
inv N99P_3 (.i(UN_3_IBUF_44P_O), .o(FECBUSY_n));
inv N60P_3 (.i(UN_3_IBUF_59P_O), .o(GTRIG));
inv N58P_3 (.i(ENWRITE1_n), .o(ENWRITE1));
inv N54P_3 (.i(UN_3_IBUF_53P_O), .o(ENWRITE3));
inv N52P_3 (.i(UN_3_IBUF_49P_O), .o(CCLR));
inv N51P_3 (.i(SYNCLR24_n), .o(SYNCLR24));
inv N45P_3 (.i(SYNCLR_n), .o(SYNCLR));
inv N94P_1 (.i(UN_1_INV_93P_O), .o(UN_1_INV_94P_O));
inv N93P_1 (.i(UN_1_CB8CLE_3P_L), .o(UN_1_INV_93P_O));
inv N101P_1 (.i(ENWRGT), .o(UN_1_AND2_102P_I1));
and2 N105P_1_8 (.i0(CGT_HIM1[7]), .o(BD2_CGT_HI[7]), .i1(ENREG2));
and2 N105P_1_7 (.i1(ENREG2), .o(BD2_CGT_HI[6]), .i0(CGT_HIM1[6]));
and2 N105P_1_6 (.i1(ENREG2), .o(BD2_CGT_HI[5]), .i0(CGT_HIM1[5]));
and2 N105P_1_5 (.i1(ENREG2), .o(BD2_CGT_HI[4]), .i0(CGT_HIM1[4]));
and2 N105P_1_4 (.i1(ENREG2), .o(BD2_CGT_HI[3]), .i0(CGT_HIM1[3]));
and2 N105P_1_3 (.i1(ENREG2), .o(BD2_CGT_HI[2]), .i0(CGT_HIM1[2]));
and2 N105P_1_2 (.i1(ENREG2), .o(BD2_CGT_HI[1]), .i0(CGT_HIM1[1]));
and2 N105P_1_1 (.i1(ENREG2), .o(BD2_CGT_HI[0]), .i0(CGT_HIM1[0]));
and2 N104P_1_8 (.i0(CGT_HI[7]), .o(BD1_CGT_HI[7]), .i1(ENREG1));
and2 N104P_1_7 (.i1(ENREG1), .o(BD1_CGT_HI[6]), .i0(CGT_HI[6]));
and2 N104P_1_6 (.i1(ENREG1), .o(BD1_CGT_HI[5]), .i0(CGT_HI[5]));
and2 N104P_1_5 (.i1(ENREG1), .o(BD1_CGT_HI[4]), .i0(CGT_HI[4]));
and2 N104P_1_4 (.i1(ENREG1), .o(BD1_CGT_HI[3]), .i0(CGT_HI[3]));
and2 N104P_1_3 (.i1(ENREG1), .o(BD1_CGT_HI[2]), .i0(CGT_HI[2]));
and2 N104P_1_2 (.i1(ENREG1), .o(BD1_CGT_HI[1]), .i0(CGT_HI[1]));
and2 N104P_1_1 (.i1(ENREG1), .o(BD1_CGT_HI[0]), .i0(CGT_HI[0]));
and2 N35P_4 (.i0(ENWRITE1), .o(UN_4_AND2_35P_O), .i1(ENWRGT));
and2 N44P_2 (.i0(SYNCLR24_GATE), .o(UN_2_AND2_1P_I1), .i1(SYNCLR24_D1));
and2 N43P_2 (.i0(SYNCLR_GATE), .o(UN_2_AND2_43P_O), .i1(SYNCLR_D1));
and2 N6P_2 (.i0(UN_2_AND2_6P_I0), .o(UN_2_AND2_6P_O), .i1(UN_2_AND2_43P_O));
and2 N1P_2 (.i0(UN_2_AND2_1P_I0), .o(UN_2_AND2_1P_O), .i1(UN_2_AND2_1P_I1));
and2 N95P_1 (.i0(UN_1_AND2_95P_I0), .o(UN_1_AND2_95P_O), .i1(UPINC));
and2 N53P_1 (.i0(ENWRITE1), .o(UN_1_AND2_50P_I0), .i1(WRFLG_MEMD15));
and2 N50P_1 (.i0(UN_1_AND2_50P_I0), .o(UN_1_AND2_50P_O), .i1(UN_1_AND2_50P_I1));
and2 N115P_1 (.i0(SYNCLR_n), .o(LOWINC), .i1(UN_1_AND2_115P_I1));
and2 N112P_1 (.i0(SYNCLR24_GATE), .o(UN_1_AND2_112P_O), .i1(SYNCLR24_D1));
and2 N103P_1 (.i0(ENWRITE1), .o(ENREG2), .i1(ENWRGT));
and2 N100P_1 (.i0(SYNCLR24_n), .o(UPINC), .i1(UN_1_AND2_100P_I1));
and2 N102P_1 (.i0(ENWRITE1), .o(ENREG1), .i1(UN_1_AND2_102P_I1));
endmodule
`uselib

module gt_counter_globals();

wire GR;
endmodule

