// module for a jumper
// MSN, created 7/27/96  
// last modified:	7/27/96   


`timescale 1ns/1ns

module JUMPER (IN, OUT); 

        input 	IN;
        output  OUT;

        assign OUT = IN; 

endmodule

