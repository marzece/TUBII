// null module for a 10-pin connector 
// MSN, created 8/27/96  
// last modified:	8/27/96   


`timescale 1ns/1ns

module IDS_C10 (PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7, PIN8, PIN9, PIN10); 

        input 	PIN1, PIN2, PIN3, PIN4, PIN5, PIN6, PIN7, PIN8, PIN9, PIN10;

endmodule

