// LED - Null model
`timescale  1ns /  1ns
module SMLED (A,B);
        inout A,B;

endmodule

